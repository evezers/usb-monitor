--
--Written by GowinSynthesis
--Product Version "V1.9.8.11 Education"
--Mon Jan 29 08:53:46 2024

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.11_Education/IDE/ipcore/PSRAM_HS_2CH/data/PSRAM_TOP.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.11_Education/IDE/ipcore/PSRAM_HS_2CH/data/psram_code.v"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
xTU5wEOwQhnARwOmXbJMNVBX8a8J0Jl3gR6Hy71JdGhRH31g5NzxR/e0wePatn2UXG/2CZ/0dPsI
m2AqcBReUlbXVHfIgdPHYCZsHvCUxivOiw7ZUchFu/lj21feqfKvZRlioTp/V7YG+l2S8Ux6QZvq
ohivAAcxSo17DViyfBB9aX251ATKXXfM2H1u/4534ZXsCnMFmdyMm2mmb4MzT0az7+660pT9ksVN
gG0nASNzHVsITHyPSQJZEOlHVGhBVhRsuP7DiZqpnmzBa4Y+65Tx4aDJnjDk19GsIEG1Zq3k+Evz
BiuCV344CuBchglVrOSuG76zJ1Bfikv7OeuX6A==

`protect encoding=(enctype="base64", line_length=76, bytes=373168)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
iusrbwm5JZxy64LticywJnHXXQX0ZNtkBfdlgz/n5yNU5BFa4SV2w2aivRSIkEPHture4fRCF1uf
9ycFoU/53VxnpVWOfMiWTtFPIS9CSyEEZSodp1I4qULeGIE42bhyxD5kShl4f5gRxPjn7D3qtI5M
UzyF9O1BUUks9fq0ZgvEzGbkwevKtWALaBEMhr+XWUkzYihl2Fx8KLLM1I+IREAxGzj8R2lbOOez
l/q3CiZyYg7P61bp84Gl4PAjg+F5U07/BuGnraDpyx4oSuPNwEBKppvE5d3lqZ8PjjqGfd9aG2JM
Doj3E8J1wco0l66lFGA30KSZxsKDob/v0DIAHPt9ekKEkmq/UoC8PeOMoXSxw1gvMMJdfoyu/w0h
mMK2YK5mLqH/BYZo47Csoq64SBthDagqkwpcWa1M3zCndfXz1+v3jlPOH6Xn8pDnwj9CsVFakF90
h3LJiMISJCqzfv257fC+HZcjKt+/SHr5pOSwKEUYAdWNNpPcqwtWoV3AZOQoMixRaFxob4k9vk6T
8UpZPNZTY+jGjMPzUsBWkPo0bDNuAEBJYmXXfNdMZlH6bLv523DLjwNCoYZ3OLYj1cYHPysWbxZd
fTlewaSPT4RjV1oNPV+kDVyyQtra8+EhT/g8PtC/y4cFfYtqkmZo/dAxsmV3z1AzZKNn1Xql8NZU
8fVQu5TbK0JWe/duz9ijOpZlpZt3J+6kx4cuHhalw3RhMPY9xwDi7BFjHSDAhEoWAwPSdEYC23gs
/rbWTd7OnguGD78kIF4pbDrIno9RaY/qvykdPIybmFd3Jui33nfDfMMPxyej97iPVQfncwYuf42g
ZQ64AoCGSiopilfDPWh5AmfRKF7F5LzRTcM9Lqvj4dNArJkRHCV4QaHk3e/cIq5lfl626f6h0y0o
gZsEao/0FT/xEWp6OesrR0pMR1lCcRTmC28xkWO/KvDUiXcyWmexGJEpvaVRK0pzkmG18AQqdMaA
QBhGdti3YVWm6usRTqvUhfQaDbbMuHu5DIr7n7bB0Ji6mLcuwjzzyfqxTj3hLRvhL4G0fJP+4ztK
zRAyB4bJXbq7Fmx8yrVueyItgnDwh58C9O1Y2izXK3mkLCOjmGZ+uugajKbXO5c6uIul448z2kdF
cCSrpIRbcyOFvbEi3zGaQbx7StndFxyaoaHpxl77qPb0j1XsxnCDl730c3DGV69RJdOcswfvaJRf
Jgq50e+1cDWEWWeDrCZBiSITxSr+UAzx7Pv2Vp0qGaKv7jGCTplu69RARL+GqqD0IZXGbHYMuWk1
ddwN92ibYNCRmIOz/0DJ8Q+mpI0mTpTbydxbTzBgWlLNrkR+jygtBAGdjxD2w605bhbs3HlqDaVO
QIrKjFYcC8EYz4+lIRIpDTeDMhY2otCAWDeLnUcW6M6NSO6Uak2NYpRAd9PwVFMWxVIL8fWdnJww
C+Ji/Cpha978EsQsUnseEIU0cQ/PQT6moi+9P6h3NjwdPnFSvLat4+PoX9mRuoBJ+Auis7uZMhNi
EYSCnwXzQUc27ntNN5arNJca6Wi5bTKBajV4HyXM5vsYBA8sf0bAEGmikKx4DPTmfSdpFdFBlZP4
IvOZI/xAnCp5uzTLvvLDw2qkN/MjkydakvuWYGaumJTnmZnfAtZgsq0otd2Swyxo4TjoWSRiFN+w
U5j+Kv8XZs4gyBVRy+y+JB25n4P/CYBXMLBW25pEc5Q0K+OtoBYk/D8+X4K2Sy+SEu9lFNx8gSFE
SI0vAzsO2nwMtOKUsuQHCZdr7oWOntbcZvy05AsFfDqD0LS2PNZGn3OvtB5mJCN1wRVCzDDIcles
bOTB6/i6afQKNpuft64KM7C78DfARiBHwG6RHuGmlMwXIe942TNPcyFSKG+Ap5BrXRo7Wmi0FZjf
OoSCwkr/0tvuyValAVqUQi9oy/d9khLemgkdsY/uV+a1Kxc4+LZgELX0ox9ngNVoLasgFD7iUyqm
kYhvvaXb4ozVUhLkmsUMmvHeqSvsX9LtqBBH1gP3wpCdD33BJZtyi+6X2i8d2+uU2wzmzESNjZEr
TwzXQwKLCCDBfY7590JLplamF/sukw1Zp0qEjEEBccjh7jU8j13FJWYnYA5Za5rldk0rBH4ylJg8
FbEzpKif4FTkZdkctDJm0US+4ZLU0SrrSk9g4oZJ/o9092RO1ZM3mYEsEwkHjO2KC+yo3tqG6Xxh
16IUbsnoZN7ifjeVDdJnl90MHadyGk7Aa221KFdAEmjrTpzJKs+SmqTAqjSqS6+Nb97RdJGljSH+
wvNTjAsNB99TcEz0iJB0Ydhnln/qZy8+PLrsbrtJ1Y29WrhTeWd1H2yF1IuWu179TT9KzX40R7gA
u6lNz2/eBiJLyklOe9Y89jtjQp9BTncNC/6F+bho+fT7AIKL9kB1gCyhfe92JIJc+H2GRef8hPqT
UaipK0yJIzc+C15NIAZMZyftD3GVklMrq3R2YZQqlm/APtAoRkFdv39Puvjyx5mzniQWObT7Beb0
a35CCOiGrCoUf4bRVqJ7rBGd4//25XweL0KlRwka9JjdnsmMExkXSccAhLhM5NrK09A2ncvCLJIZ
/fz7hKnizN0X2M++b/CYKCl7c8AAu/Xf5FSd0Gb0rEnQO7koa+A+CSlcV/mPrWRr5HbwfVhVrl/r
GUP+9qhCu2KcOn2/zc6esMyxDFrwbHnCHSob79P4J1OJx1HpaXhWNOKsMoLik8grY2k01Mi1fpe5
A9Tdw/dUSCCKp7JmABMBPwSxSBR4q3Am9Z4I9A9tRzRc/kvXvvH5cyee33LJh68a1Ay6n+nIH4Ps
9nnVBHkXGP88vAWeHdfk1RqQok47GPYdU8YfNpGB2wUtHqCO8qXkuN6x3w3xKRJVQlbiJpE0EBqO
vAfR8hIGOPwBwIDhvJcUc3IVFKkvVx2nl/W5J8h6seTgne0ZApJVO79lmvFLr4EJc0Sk8WtnXiDA
4r9AipAyIrffCOlp2s7rRyGEWFa2WKl8sasp8aBG/ZfQAUrss+6/w+LF8dgNgT21k1hWB1pVrqAi
LXM7fVwOAezNsWVMjUmZO6CJQ1Xz5gw8f9OR0pQYNZJ7Ma3XcR7lHTwiwN2k7FtVIJzl2mom7eI5
87mDvMYiYM8koPAOm5h1W0aS8f/L6fsR/he1+jEwkeeswjSTA00zPPBd0KZbbasq0I51M9rFJfae
DQEUqnU0NXJNkZUYgZXpfEJXWBHRLsxWPFT062w9Pi+IK+1BKGIfiRp5ufqzjmXHoJjmZ34R1tAN
p0NoyB4lkhzWDt6t4F4W85CiMXZqXzejexHgaa1gCKtd6bpkxxiTYegA1MYcimQ93mx083n3rHpl
1WBtkT4ntZ+zLcf1umyCI4Zh15vbR3O+qC1ZVShe6g2KKkJduHYsWNGaEnHa6GJ7G2cKWaD42QEb
EqtE7z2H0WEp/RYZvnTDWDcNOcJ6lhIRL9T0G9Fs7sDlSWYAMSd5N7/RBozOxrSd/Msz4KseYIno
ndUcdcsB0AOja8HoHF/CvGcF/+5U6ROoN+V5O/eFC4sS1qmoN93N5IfkJ9xETg57tR9zUAYiYHSd
Mz6+vI1pqewtaLR4SK8me0PTo3dZl4sp0xHhpV54KndgCm8IKdvT+Fz50PLnKV1RJQiSTNTPHdu3
MzSReSncyBXfmTXmJYTCUb89wVttIppIqDnYSZnzkiiwGDvMt3VgPsIzgxJqehQJBA6bc/ntxZly
HEUrHeuOFIDKvHmkdcjh+P2xlZMREN4y4yk1G6oJf2x4+jzRhe6wDJ5Zc5dG01fAExboYPWrIeuM
71FlxxQn/FwxOO8CGn6iCzLBw7uqXvxFqIpwdXKdz7A+bJG7SAqie9CSjRqGIs6kuvOizQN8V2W2
C/3Dxo1681C+pfrU6EvbuFSX3IiJiIGpcwLMN6QwViMN+7sgbw7ZfpILNYObNC9buj3XmSKJ+ug7
AYfb+0qN0Q/+8P3oy8VpSzUzelpz6wYJ5ViMnyhs2hUC0fCF2grQoL8p7fYOL3ne9UMHz+S1/bE6
3ncW9a+nb12/lVxPTdkZb2YwdZquWbOm8jmnz2V0ZyidB+OZA/cmWrMQAgxAT/Qpx64YnlOP3ybl
eXUnPWhUpxHgf0Nb18LE/BZjY8udxaoa4VNCAJ//N4R/Lo3IQjRGKzzmQdHKxpGa7XWEBdydO8mJ
VSuOUX8Vh4ah6U5QTcZUPMZtn8Wn6FIRCV72KTBE6adLFxavu610bIOmXnIXtqEh77wCwa8P94lW
vLUfDNX3abTCo/jaehH0MgUPjrRccLUmdC09HeCIuL63EKKeCKhfuv7l8hoRZgJl3weoPCF3moeX
fp1Iq2WjCQ+MfG4yvwrHjgip/xN3UfGrp3fW0FQ3sgx2XojJp7vv4zGHw800/4nAckSRLLQ1cdZT
kn151T08CMvQVXzz8uWpS4/z+kR4ympbXo1akaJ4YC5NVmQ/uC4sz8D2v+lrODGbYTR9yy5rkFz3
RpXL8cCMqxselJGokcO0Xg/ortUxMQEyWWQUn5SubJ7I1jYVZlns5NkllvQ6SHACwo2UqkrufWoF
KfvWtegUf9SDQ/O358hv5hIQPdFiQpKaq8Ao6YGtv4g5uEg0UJ9vwiGYh2oBdfCk6knmt+vkxuJv
8RdBxAr9OByvluz7Ly8YWgINTeZpaMTkjTPjNFagaeosB8/chvS2R4HrW5GW7dfQGhI7ZBSGy6/I
Iob8T1+i29odwE1ZSWajna5lZ/Bf8XoX/qYmhe6FDXUrCtKpvu654/xSqOwyjMLmsX9WyIcjUOgZ
iSuffQUnZMOb88bXAr9iq4Fdqwn5iaxZMirBdlHhlTX8dNJb3uzmXQwquC7NmoB5Fvl9WjQod/ZQ
7g4ZABjnthCt+VgoZKhkoWl820fP78IVhqYtOFVyWwFJGIIePT5/oai+3c1tM72blL3GXG4D5M/c
b7TIpxx0tYZ8zs9WU1qsWy3zZp3OaggVPmasWvVE2Y8148HtDVyXCn6sMqqtaNnk9w57570X4zKO
0hQRsciMffLWH9bTzBon9XIHyLHMj9wjxuFwdP2xEA77PpOGlzkIwFQoWHaaGTMnN7euwt8mAZo7
lujG+fL/Dj+3e15N6mynlJyhCON6vf8VXzW/2Z02Q/LkImusUAMG4VEitlGEeCtNoXsMhQMejj6Q
hEtqcu7bppk8M+hHSkuHcIL64VTXTv4VNDfnSQJKhO4DR562+Xx7DPikgwOdV2lsZdurY1dopqOi
IhzsNy3t5OQBYYuV+Z7ow2lNDfpmdwG7hpdEOO+ksCc/gkECXy7nDPTUtZNQ93KGcpBn8TH4DRXN
17KDXEJ9JixZZ67eUbbgjDCDJOnNTghm7WM8zu2sLRchWW9DTG5FAhDBSpH6M27irPFmCYIUA6Sv
mNusajCL73PW4XjGG0yMrryaPIi0gSM1R5uVGBBvGJcRlGJ9UYUqllpDZ0pmakGNvmev1ZlINR9b
Exc5DJGBZVsnh/zmRk+6vzC35PJEV0O47dK9P10p9R9GhvyyIcVwIEi7ofYm81pd9hQLPug4ifa5
SrYD0nS6C0t8heZP+RxvdOn2okk7vrE9exOpTFwkL3f4AqJ/RZ8eE2/1XkxkHveqdg8ac/CB2eag
lxJjxivhdGTpLHdCTeKf5nowcgfMWWTO+4gpZqz5eZ0LFCYNfiLQ36met1vnIXqVMztW3Ea6JA9U
6NRs/N6IwRmBgxQhw1H+OYAbFFwaHMj9hmHr0kv2oXiFULOZnIwgkjLxCUeZb7mUbnIjMlaJiqUM
P1+BfIwPm8/mqIwaDDREWt4uzfzyfKAqCPBuUwuPnt7EXOSPVz77wIoyJn0BVosWnWdz3KLih/3G
W971Z6zt1LY6hPkRQFjFP096WjVWasduvJ234WMQmIufSWh6IWZYLct4vMHBSZcyjLWN9mmH7DoL
7zFATjv68bMZC4hKSfIZsijf0m76jaHsV1l7fTVuWanBfBjN1dVGH4Y7+/eNUhBzY45WrlD2tk/K
S+BFcibaIvZw3Zl5vwuvyPy7K2P1IaenDUM6qmWd2Z1mkc5wVMY+vGzDbsBXOXMp9dqIq9/SY3dH
zM2q/YWLoBty2DVGLtDEZI/zlsmZ1gXsHI8/kjPNTZhLgataaAIqxyrzW3Ff/fv4Up4LM8zoEWBY
Vjn0z5QFWXU8i/9bzzkybvBfeH5dH5b58NPGI7Zdw9kTAoESJPOpjDLLqxIVH6BMUuDDfZSDgXYJ
Lhz/xwVSe0p31UMHKHxpiQEnyALLXzqBLuNa9FHDv3AU/kBy8IFTHmoAUJ4ZTnIFYjLRxR1DB+EJ
Khwul//NjXv1Go3pD7jDWUX/0JgZEzC+wPPaPprCMjwsnHXpPdDyknd4RBkghhu5niKxbRTGgM9V
BFFCLoGMCsrbBoIOMWcGpPDLBOvNvhr2Ef4dvUxiPF3ZisjjXiQRptD0++nJ3gr9t5Y8Nae/s8hJ
zNmOrDrksnIcYcRToCngTRsHo7Osws8Ql0jk17jMx+dwp3q4M8fBbS7Wys82ohcgbE/8vfs4Br6V
2e186LTm+Mz0Yuwr0JwGcU2/h3ysVBD06mhNN53ifpmN/qLmpe/jYfcP/JcaAMb4qNNYCquieru9
vMkFM17VPV17AXeNt0DkH91Hqvq1IY4kMCtLNRc5h2Gz64uR8/JDL2Xi51/9iGZTKC/HbgCdtBs0
8k+3NndhzDCLJ9oSRTsRho5wBZ//5aJn6lQb3n516LqZpxVGBWdLRUzWLlfQg03afHaxhKsHXSAa
xSvQxt6iM/HzvHD/tfLgDGxewjvXEVenjWRy3NuH+L8lRBXVJZB0pipCqp5ThP+dlnMkabRtUhzQ
f9SVChFky9020jp3T8k7SbTDaVwqkJXaEhEBh2ndLU8THYlkJiC6hhRMzZxQzQkHHqZAkEz+9kCZ
2N0lfwiWhxfk5UQQd1aVubpGnnhCeuFypZm2BoBQlOd4YKyGdEGBNzkuJ8lK/lZ90VyHM7D/ZPT7
KJqSpww6xlWAe5XVEuQAmWdeV236gOA3vMh9jJce+PVN8fbT5qTCNgT/hcMbVoS1llMJ5DaoM8Z5
6lwUkoODhZh81I/FOXCtcR9C60QLgISOrETKBY3rUb7n+U+7gfYh7spPEnondTGCUC/KR5a1lRx1
pbhELV9ebpr9zSWivhiUoI+tmVVKfWQGikRBHz2YirpEJHqgqCf4uQTEg31q9laUrqQE8Qz09jgK
szEsughcqyriCArC73+dlyulB3zgzfnz4BTqLvOAsJ2dkSSVsR7P0URnw7oqkXsXalAddI4xkUUd
hW6plgBXqFJyYFl0vAgEKj1OfBbvBPgcJMwsr8bfAlFYCZHvJAGfEVcv4tV/aGrrUPJIsmxxqBi8
9rYaZ3Js5vylDtMKP5wdDGzRPerRlhwDzEgjF8KCoEV6w/IS19U1GgyfPx32H7YibXVapqpxYge1
FjtYc3OaHBKf1FqB5TU8SXYVd1wPgpgUVGugMLRaaDyWla47SlBBmhU06KaAoB6UGCX5u8pyEopm
F7szEFC3O9rh210tEVr2aLgo/3eGZ18fmolO5qFoAr10oHXyUVNiFVFSKEI7fNzMSMGdljaM+o5x
eBpK1jnW6m5jFl5CiU0xlb1REkNtIDM7N57CBwKuAZJ++3N9Vb0jRhVzLoSIqh17CeNMneBWbDbv
6plw0x/gaWQz07se5BWo/tYymFFsLhSjk7kXp/YN5h23pdASmeoo1RR+I7QPXsMO+lvMSu26rWVY
BXf5+8Qf7zexAgh7HCuFfFPI5lDOSfeKZBx+x5V5lnRfQftAAx5WvzbeiXPhdQWCawcOBKR8TLds
qwg4H60OHKErAoiohy5pd+Xt9innFUa3r0mVraN7TJXmz5kLFKNK93+Sfds1w1yrRr1QkKqzmmOI
n+GG1Rtt8jJiDQd6hSitnAT0Ea1xj3FYCb/sOgq2qfGlo0wZdqHLFflCV9pqAoAnPIK9fy42SgZ+
4LC3b23dSe66cnk4h4PlhW1KqZUKK7wRhwGdcHugq1J2tdQrrZmpDNSd+vSq8d+z8UHrXaf2cxo2
5mmga3YHIsALxP6cQdVSpHcDnFn6jF4OJeTj8lWEyebeht8HmhXgmqclRxGjwd3xY5VQQatPXAHg
Zd7CcI0s77+aqCC5WtlQ/xv/qiDlz7Wu7Shr5wywG7DbSIdjja2Wyd8cUGil9RNN08MVVYxC0gC+
7VgVQUAaKv+QpseeVzexHI2zKD1jcah7FP5XhNs/jCFqieWywcRHCDfNEGbFyFOlsI+zLEm4VngF
BxPdqSDSnCzBEX3serZmvrZ2aI5oRbZ3GsF5cShsWZylDDORti8JEIkCBEGC1vteqvV5DYPqIZ/k
fcZ9LHSa2V7f/Q+K30suURiXJZwedN1X1lQ0N/x6xx3LOSQcjAV7XIJHcUDe1A7iopB7mrZj51a4
NLb0lekroRHUUDwwc6mvzB0zPTvVyo1MVnh9J6UasRHtqZsFOmYBp0agF3YGwqCI0eUXhH6acEA1
WMDi6leNUdiPTIFeNGm/1iVxDyanu1/4ugPGBhKy4jzLNjquDezN5MvxftYsNTNLAxU1pbJC4+Jd
cEcaWuPCO/CmPdUzKGKm1bJhw1lqq7ZI4gEX0V9VTRzupZFUts8ZEAUh8HDo4ogEA4O5MCXYS+bd
pm7Bs7Timzst3qQZrxK9Si0+4taNAqGBriplx1U7TaldZ3/8OX77Owl45a7dZycP3SQo2vrj1bHE
pd8Kp1TeHHUFphyF+H/Gkkh7o0qBJyZESEe7+p8jjkTHCf2UhVZGnkWU63yQ8nFuqYtEd4Y4qfuT
3JertVbZ5aH4f2R357XBGzh7GgxcpAsDtFxuo9I0IlDzwyXHVGkX86Fis8ygG+1ne8EC0U4jo6tR
ptNFsbE7puxF21vinKUu87Fo9FyEx/WEeNrzNHg71UUEo9Gxr9slvf7IlyLoIxC/CbmqaOji6dZb
IqlZYDHLYGAlhWMC2gt9R9hRBRDPzCYIuQZ3JAFr8UqowrXmkAd6vVfSz2SA+eLwEcfafrLqwZ7K
gE62iusDXo8rTbPaGSiVc125IATGMqhLZ2HLFjX4kb/wdLl57QxNwXO1Snu+0s/b/I5tyPaLBsYb
+pDmypX74/UHmTa0aDZr7B4o6eAGIzWnq82IeGgLxQHCJPZNXPPtaxvcb8803/LHdK9ybcA7zHsK
VQ1JHfaKKVFxD+oj+Q9bHPL4k3COJsfldR/Dzh2bLii9rNe+m2kdSGqguhpau1bTlQeZ7MEUJgRA
wEoPhmoY1mWBdWFUkYEcKUlOn7gx/SqJydRQ/sunfsKSfdrbqxfK0BePkNvJRyy3pm+z9wB04+ZU
wUsMfMSMhlyh+8y2pHLZlCc2hKrhrbum/TQL0QWF/x62C6YfO8/TlcFxJ77Auxxj8+Qg1Lx+79w9
fR693Lq2vA/43JKtVaSPy6cXJWjRRP6alqU1O8C2YeQpSuSq/V9cpb5SoJutkvIyy7V0DMWRfm1u
xE1JclEEV5zwl70t/94tprYY7DW0K7Y6PlcEBKxq9d3gtVP0yTzWE2Sq4n6EeEO+C7Px/JfCUpsz
0GEja/N+3/V2J8M/k5d3O6zJxU8/7/p4BUk4lDacNrMsTyqr65xuuGhSvmaWEeNoI1aVV1iWjVLu
qTLKlA06uGIDfzh+emi4VXTx+dCwFygI0UFuXz4xb2hQRt+tivBop9UOwEcUk1yKhOUc3mtIvFgA
OXdSCEdvUOQD5D4soTMTem7rSWObf8ER1EU6KZULkk0bMDfsjEEj/E6EL+w+047n2xJ+x0adNPXl
x7xys2rFoCKnQL05RCBp4nKIjaa6zW/YAw/wtXVa5YmUe5SHYetJmxHIbDLbJzM4Pwy9vlPo4+EX
j6LfmjpDFCfq72zDln5/086iwGIut/+XSbIUzqpfUaDP9IasRBwrZGrLCLLUTrWJK0GcyeKnAj4b
anySZMwhrX2KvDNjzE7sx/436N+cZAD5Lavd7IAwzDaQEv3bWrlKgdjpbE59rHcYqgVHUz+BOki4
FDWpMPqG75kGG/JwNza3TCYaZ8++BjZA2IdJaCiEsSRxOxGvkMPFlGdsH6ppsCBtByfJRbvhy7xh
PrXDLgNDTnKOPwA3Gicg6gQ+3j3KPsWmllbxMkVM+AoZXjuVmhNhIEg3PSwqle684dLzv2JPEN7g
wZqaJxwB5gJoF+oMLTcDb3dyEuLYJZkxynuO95OShQqheWawKKIGzOp3yKFK+uldo+3qh2wgC2pr
al6IORNH1+TlfMZ3/A3RKkwmIWelkpdLmXV33q1I3TVFIWf/wLJsyw9mcAFAldnqcfyFx+qcLUKS
RlxEs8wD01ITumkj1BhvvRaY6iCwTXKCfitJoW5l+nljQAyT+NWZoRZYYTFFj8+8Ht9Nuug87bOC
ubZokKTOo8JtuZW6VCbbQi4AO8nQ2oHyVV7caZmGemdIJ0/ssFRf0oKV5uKMnJlEjGUKk08cTVXU
xB4nj5cpyyM/gSsmDBcmtCrIKNBlju3oBcMUWqm17Y0PUGTznygZDWi0cUbrUoJYVIU+GmkM467c
bTUwo+4KGeKS9k0nB7rsa9/YrYRqntwBTad1QxBHJ4QHAcQhqOyGL/HgGfgmKaiDPy+O/cMSskVa
UcO0mrkEpfHeTkBrqXfWqxQlqBRrz0mmVEco/vbAMR3Unw2F1xv7mvwBBQ3A9fTB0/CewqXCUhjD
J4SJ4PQH7IK4OuGQS1VL+kK3g4EpgvsXQpmzy8zYUViM+fK9ph4EBdWyjOfe/ZsqTYWQrwzHwbQW
1r+xhRJpQNqMdyyZ3sUSZUFw4VnYOAeCR7y6eUIS9hlz8T2yU98PwwluapR1fRFGUFhpXCIqj2qf
5mdYy5AUEWqcZMZjr+b7VNfGOvk4HJuUC6n6cNy1LQvIY1/UOyJyWI09zWBmYVM3sxZmeaV6TsMc
vWUf9MJrggMuO5yfZQbzyIww4BfoxW7iN9P7SqzelLgTnHbxjzaFqu+2u+IYECWgZNUIcTf5vgcF
BPpspDa0YIJ2tYw3OxKK6eZSgeuf0URo4ChtyugUQN5I6a+v/3JRk4bCXkyBhzIRVaSQprlejTtg
Tox+vRfDiNOhDXuY+cCrI3u545mZiCtnWdScrHwlRQmpXDP0LT+kVhXiE7ASIyH+ECzF+KXsOivT
mNAJxawv4rxezYBjWIRNdDI8cJRH9Zs5LNUbk1UQ5CkoXt50IY2vax+ftFE1SuCiHKiWitE1BBxf
MU8I1KLBngZXqkybrelntKDz7Febs1h2XYKDdKcsFExoRfxG65pyZQosA9rEWJH4ejB7eBJHv/7w
/OLGm6KGH+m4WkDKWcRhYv0dmbOHRB1/oRo8WEbAVRSV+H/Weq8OtG9GUFpz60s0PcAEJVNKEjEq
qpVDJY0EI5NJBrfA4H2i/Psy5paTJFrVPOUR3C7UDfsN518lZmSgkOg5mJwFC5pXkjRHj1L77bMW
MnU1rVktZ4QKHboZMsrHoiE6v//lYbPaQFVDilV5zzv5iU3g4G+70tnRQFbhTLjk9GsQhoc13HbR
mDf1nuS2vgbyw42+MCFBXYS8I0NY+1It1D3MgWWNwh30ui69r6zsmwDnPiBLH0Wql8QvabmS+wQp
vvJeWiNgg+6LEH8EVS3og4lZ5MjSDJl6QDfHf5QB0rcutKS5OxdJRcnC6eZj16piVoKHmx13snFH
N+6nRKxuMP0zhMtMMQwzEjkssYUQFBI5wpG8YYFQNSJ4yANywbnclIo0PAmQjhcH+7fu6u4yqLX8
zB1JiyNxbKiotgIeGbL+SEmpG9seje61bIWSUi5GR+zbQBkxeDGW3B2FOuLkoB/kSzhQd7j2arT+
i0oRtJiWDEAb/DFZKaNLNagWBoHgB9Zb7MexLsm437pMUiY7WVbUHpkafGkhA4JhixmcHVtSLUXJ
XJ50NFmYdYEM+z7sEWok0wRpBBw6yB8zD3XkuZ/ChgvtfOAqJEEwd4v5BiyTdlmD1pvLjE/f+/nu
zqVsJ6DMmwhHpcOZydv+M4xus8WN85rvULgeH982KRjHlunX9auaMMoJZLy5tDNYf51/zBvED7bD
t52rG/Ofr9T7Blq/h0098kAEyB6N9vWUHEuT7pI0yh837X/Fb1oKfXT/OehjE2M26Pt1XGpQebi4
z2e6gp4jShy4Lbkqr+oY5dM240kzklYuroT7ee8JG9WZEp6ZKA4rdYyKPk2SVhYuyKWwsMHWQwsf
nStPmSiy6L09r7cpQxxfiHQGdigD+rU2zFKRNzQphi2yzh2stLcky5YBoM9wlLg641XSeekVDmZY
yMuwHALSlFoJZDoQl3h/DhHajRqNHeBe3i7D90GL7Fk8jnlYNmWCD2jzQu9FCDA2Pdn0VTJTyFtr
sV7eL3tiY5PSzgDU9sfDKH/LYgZBxBGxh5N13WRlPstak3K9Ha6/faRCsmFAiuHHTuqBww6e+Z5r
vy3qR0xy/gteZD035BmoyaWJkK/lEZAIi006DeRnAY1XiClbUmMCHBJKPFKRiij5X8P28UimkfCo
1H0hukshSgDce+H59gkgBcP4nlTe4G4pa/wALCVjjC+CnSnkV0lB1hfu1S+SFbSZsIoa2CNrKtLR
37ZVdA40/1Npsh3GoS5DzK4zy0hHOCZ9IoGdWNCV77l2GAaCw223vtGmuMgjDrk9f6S7hCqfAwZ4
U7ORLHvV+bOzSMVl/1AMMx2qtoqzEgipMB8okZc9DjhfVv8rvu7A3JxqC7QGKUYod/G+OCbSW+jK
oK/mPdQpGuCPhe+XamX6Z4bzhKduJkh0/YS2jrhte0KXlDXE1vCbtEmolpj5R1nvVp3q8I4hkOCh
LSTnozCSeImHMU27osiBwNzOl+K3qmaY7iKpbfx/48k1oVwxILGc/+vDrdcA0wPybnBqDJ/j343z
gK1y3NfurkfIS/8YDstgY/N/6ZZBjeo1Ti1k+nerz9mYdZx0NAAnselGtvJ/R4AVa4ANVznJnUF0
Xp7omYmLI9f56dPmxXNho3lDHc9kd3zpj4Pf9yZbTsrJL1Dw1wmKD5BUUoE7vfK8CHgO3Zo1je5I
sAtZHDDIL2AvgfSjbTyouQU9mQ7eNrjqJjKhF34dPLxa0XSNpJqpthli7uvVe6oBKwxv8qWbGkXt
OX1y8BH0SqueQbCMDhQ2iktZW54eAEeb2wlKS5j1lVD2l7Yv3T3izxF0jbirQTCZ649oSjhqOYRn
J4SPNVS0CRx1ZkVKi0gjdBIlWZG5WyXI0RHd2zGfST0NsBvQL2TGELU/GcBJ087jP91ggK3FsUvI
+5MCyRFLAgwR6BsOYV/rayEib2QULMNu10xWSyTBYQ9j5su1Sj4ba3GU5EqfQunS5tulA0iKgDbG
YO1WQoBCQXHS92UrM5ozcnOVn9UNeE5+wD0i3YJgfmxxnEdyEQBwHQeFExCZ9f9pHgzVi5AeQ1Ui
p4JDiVJmzVg2BTnr/JNLizu8Iyl36xTBGnqR7ZMFbrstyZL9DIp8A5ITz2iR/aUYqkwniigryUHE
wZNxR9oWtAB+ylwXJVKXZd37rsfSXw3p6/8ZXzzmhoPqWnDQp/2dDFHN0Nd0rUwzDf26BZpG9ibi
iNaoMOZmPmzP9z0oJTe9tuAI9iqNAJnVJrhNbk3B7reCXA1ktdxBUfpRCNL03Yw4HamS0OdkiI/0
phS/IDSnzJZUZ3UKgdV5iCEmaVu9loQ0GDcj70HNrQpS5zuBA7CsZ6gE3FuCWhWeWH39ZL8YzRq8
8pYwQVDImE0W27eXYKQTxhWdvFaIEIJYypQcBc0gt2H2tOlgmKeJ4Unfhk+2Ia4ZCUhkr6mgJlFa
udHnXd88M3LyFAp0/yzQ9jJsyxgBixXtrfyHeH5YYLAOB/xzeuNM+pwyJdbRTXRkEKY8W1l0DtpJ
EY0aECqjF5S9i8Jct5RqLRwafi/+sjxBXbkmqcd8tY6+ZwenTl7oJbkOjE81p+aXENEhpkG9p371
H/3bbQKOUv+alkiHkoU4+FtnJF2uowqptycSJXISp2YKcmM/zgbnelhZV/scvbTYkelDKDlEWlyH
y+vbfAdUzW4F5C1PKHSkpTtRhaRdf4JcC2Hcl2ON2RovPVa8BJUtpoIfMILisahJcQtgQ8AGOyao
Dl1tVXDDBtLizRyZIYQpWmzAO7I97qo+wmFxzcNGefNJ9RqtGHOZ+zA7MIo5Q19eHxUZxK7TFUxK
fv9gBkbhM4zafQAB5epiUyMG9oAN8v5DvtVDdM6CM5wlju6Pc6YYVFIuJymM2xRnSglB5+4kjyhV
DHWghh6N1jiWNiCW0KoYP84t793J3ZVat5e408iJooX/DtZBZdM9MnwyYlmAm3lYccdU6DpzAYNx
unVrHxPf/kCapdCLgOaNeSjMFUHaX3tLxI9TbdzPq6NZ7iq2jhtEVkwkKjyRs/A6uYQx4hK5Eftn
/RJuwShbYI95AQQwI1UV+eVak7iBfbji1ajvM6GU9H8a4s2ZN/UK/DiM5RzaMNT3JXKJaayW0sGX
Ab6e4Xdezi2w5fZyqDh+HSBsAuxRXJSPprRDPaGTo2/BzxyaRtuQpyi6n7ZXzK6ICDdUE7Giwpx5
6w/4xvYBbi94LACkVG4pjcnewvGlp5fR2f+wPUeFjYX2UfO+fLKQ/vpAQGJ99LFYmCkj7U0sV0e1
MpgJ5U44xpf7dWHwGb49csHnX+imzsbwzqQu34QhBcyzFQMDifaQ3qlkH0reHSLKDdXkDdMS189C
7LnnpDWXxEeAlS7mGl4E0qCTrTeXAlDKwL/ZxYAa7Xt+8LLMZixEzGy0jzlmg8mvWuOQbeN/2I6G
/+i2jhHgoQf1y0T6mJtP2ZO3EDdOLZDoRlzKplRgA0jYaevsmtZBmSgkmAOmoN88Cerbe4lw2IBX
BVECe+qxaoVa5Tx4HE7loGgF9m/rViFz+BloXt9EtmGCa/+j/O0Xbg1v/Gde6Kg8aU/r7EkCcQGB
1ZCDoWZvdxLY8URyYKEqkeJkXBRPSMgWppSuayXHgd7dOtGZUPOs7Fhin32okDfts01cY+Iw/KDB
uNc3cRPnhyACRxXyNAXalMw9oeufLiHWf8KVjTsGr4gIJZWL4K9FhvUXyOWpqeJvPf1UNZdSfS+F
upTBqJ7hLjtjHgRZuYm5iiy3VFdeVmE+7VxzKfhhe+TSzEclh8ACbHyjtsu34sqnhIsuCHtSzwrh
ipFiCH6sJIAmuK73sTkyVvtMflK2rT5xLqFu3J3RhX1xCq4DL/NU9tLwXlQ75wmZ7Xpa6ASFcBBL
FllJsiBI/LqkMd5T8fRQS3o1HnNa6TO4OOrIA7TbRF2KIRmFHuAkYMXEtPS5DJHGeRKbU07G5rvL
RRyJ/HuMpfnZRpA/f/aCUJR6tgvXdOfiCGqQKBp/8CZbMz20iPmzL33akIaidyG911kbtam93Flq
ZgQpC+/JsQ8jGdPpiwVIG2133ZmXbjaOXBfeFth++WHVvYrju7XNNsoYDgWjdN+ibfC7AHgNpPHL
9mHAc93l2PmKLI4cBmJRL0m/SNmIAePnEkm0kOGB/sJ/W2gStofuo4E+u24ZO/Z66u26x/UYYUXF
XbmndTT0Zn72p+z/5TW6kRDHOh1920fVAksCBJESr/rsmbR0S6T2jdik2f5jdWV7T+P/qYvZF0n9
P6gpbzuFk5vUc+a7cjhJD2mgUubR8CcXgP9zpp5OIR5/KKGzyEaw0uskgFO5/C4MJtZNsUd+WOjy
CkOsvUDWG7pp30ex2GKB1HZyRiOOn5tlarM3+yFZ9sf3Depi2GrXSVOhiB1d0lhfgAQ5lm9kpy/k
KlEYFGxDvCOsAyYetz+NVCxIN3MJUQeVH2nC+TcGrN1gtd6YNq8XdT44Xa2QpEUlvRFzxLsUyQqN
K9T9t4RETOerqOTPSloDepikhUV/stFm3xU/tYffmMT/4KbIvMzf3mxQqFUp4mMR6yMByBabWPaV
v34Kb7+20b+oliPlvPdy103/GyeifYN+ley3T0dBHaX1tdM9CMIFTQpDlld26zUQ/qlKZpRcSgi+
XxkcpHaPo7KnUMExJq0fuG9b5hMFfkbDpmsZfutdTDe/BWkCbxQgVsL1I7cx2rI4GR7O3Whn9J5D
c/Ytm4cw6VXPKF9Gn2xj3n+Bnz+aex0IK5MIs0IxVVMuPcJelgi9JyuGA2Y7Tjqz3VFLYHU/ArOZ
WZYRluPj46v8s+NOdA1tB2Cm2wnht3M0iIjMPt3hBYMhZN5ZjhKB3EMOFmhRk9N34k0nBxr5BeKe
nrzp2B/LZXLwam8xwybm4gvnsQFAwt24gZyYeZUziBlcP+JD53irwQfg0322I802Qaf/SUiI6bSS
UPvcDNTkb3TEEMM1xa7MFQVy2rYUFrhj48XBgFrOFfNmhKxhn8BUT/qYG3vEnnnnFylWiMp318Cf
jMjFD+g3wGyKlY99mIZR6sAD10LQR6K1ifsk1eXUUp73RwQMzvycdG23wNxhYvXu8M+u/namiRZu
w0qe2UXDE4L2LItrin7JkRTG2zZirTHK5y3xMlbGRntwEPJa6UnjySzV203ZNwR6Cw6nnJ2kCsvs
bB+qMjJ4u+HYdCf2yhl6rSFFg9ht1AfDa4IwspbZ2YHdORysgu/GK4MmkqjPRDM2UoeJnsGXQ/05
po9MqA9dkPRLEeaivD9nb0fw94vkVoKUx36zrTv+1cQ/aykWuctZJQdCM369uHTyI+jKLmUPbXZ1
nPC/bAIH532PI+/9hpnVJ+Uj+rCvPeYAYv0/y4Gyt4qNhssitnheOfGi9Ba1gXNomrbDD6fjsmT3
Jd77+jDHzrbuYdK/5rjlWQf8Kk/o8Hgkmm/j4a5NbSnZM2ao8SBOeO57T7zC0LPudYP45IM6NSU9
Nm1NG/fVFz852DMNveUPV8sLpQJlrdkwZgk1tbkJjFjlTJqO2FxysoQxnkIvRJEAhEOOKcekxrhj
pvTBXY5HLn8cnJGnuvxQj6diK+eI1DDOQKNZ8zSPS3C9PYzYADUOgFvh0z3/uKuhH1qJSb0LReBK
97JRGn5oAC3W3I/CKlggb8xqtJ6wMG12fQoG/0G1RkoIfpE6tzHMt7jsdxAvYFErHXKf8h+Tu4uc
bLpLEGweBcEm2LJfj1zkv4v1GkK25Dgge5VVhd4mG9+qxRbCteXRZAEBLmeRPAB5WKTAzvbb/wgV
LDja5bbzjnGS28nE/fkCl5lTvhV2QXv1VJKLBeSX4v9/FNVhhseuLvlI9NeoxeGzzybq+jNKe+JK
TC15YwjMSqxFF7cxaBwrCAvaXumw2ZcZguolUlcTarioLwob/Y7NrJNOttUi34SLvm+ZP3+EOBYh
j4KrrW7xsNIePqKM5lTOjIt+cmgImZrwu5hmcpn7YdYedgkWEFyFXOR1dGRT7rf4nwkNR1S+vVSH
LNYTH6VbF2tMcXs7hpr5XRaMiQSk/oMA+FStxkbaFml2da3aOiWkJr6teEEPOuIQnIYGjYF/ME70
svhlLZrfajKsC3l3pozEvC/n3U20pBgdW9ToRkmav1qXES1I8Cvv8mpQfwlNjMPiWUR6jho2xt/O
vU7QlTxGJCZEXeUPSSFs6MGoE3EdnD8Y7JcRzQVdGla9n2QnM/b5f+Sn3jkZhH4SYtYRW9Q1vcKX
FOukJeM1Z7+lMEsKvrTIQdZIbHwchEz5FSTf3NdZ3USV7/zdL3jleWWLXmfiRNRfvnyK75igaEYv
j2pL9RJplSHtT5IT0aZ/UvepuCdycsIdR+y3dV+fIPeCOEMJMJHAuS2oORVgEvwU5iYxgZRJS8Iv
AjQazkU8PwH3tWbuj5FJCz2jfNqlulrkXOBHb6okcV6V45JtAfrp8JiChtrY1vkAkDOCydXimOiA
xP2qE2bvl28MikgRyC0Ik3VOH63FWG3ZrEPupnTmOKBcLiePahtbwRD+E8N0Q/z/R4SjwaAwz1fh
1A8Ak6GmM/arXJP1RFdlbvRw4b3FFhMRtLTmrr2RjEuTd4Qn8ufVbRhhfY1i3/da3Q7hczKND5TC
H87X2JtHz3Dtvlc49A0WHVDifK3gqOkLSe2AyV88+8LfKgWARk3AXqXRid1jrhSEr41oD/9uvPjG
eXbxvhgB+IQ9RVXEvdTRqmvAMVHXxucH31MGYEaSAUG8s5qldcefAy7egk65/U2a+9nsm4r9eY3b
MkitSePhse0OxsV5Jn32jThaPiDjs3dyvGe8/0DnOJPJ0syTaCXxb/cNf2N2mWkHkRl2gSovKhLY
No3DZU6BB/Pd+mbw0rxQPEgXfh8xbI9mkFQgazYH8MOxy2SlK82xUHjKGa+VV/jtCwsyzeeEahRv
S6BEGMpJm+cRAP39OZFSSTrXBNfgftIMP2n7O8dsvMTAWIreQEEkYKH5oPssu2/RCLg4RDQMOj1g
M/smmFdhiB43IXAtYD3y0jQ0eY+Wc7Osn72ubGyCop1kCeooIfV189sS4cxi7YNg0SOhwqJVmN6R
xHsRPMu2snaRwiYzuEnJcxH/00AVW2B3F6J95VlFsRT45hk0/QvFu1BKx6GUym7bVMPkmbyR8xaV
tXRSs8xyoVT7USlSGco2TjItJHJYjV+gG7mwU5hsQn78rU/s5aBipQ5/JvRKPZGBLa8e9cLfjJjJ
kLXUz4Emk76nFbAdIXQI4nnvRg0FA73dyYLfjzhGYgcLPr55QiXGrXVyaztZdK4pvmVF7JmHGCdM
33R+Ry/6b63Txh4rbe94UcHDMuDKb2jtk8tIQDq1/RLI7sEAv141JLo8dgNBY+t2fvel+Sta/AE1
WVwNnQpnIY/IJDpBs/0zg66zccBDL9+1RtMLmLFOhtZzJTcLV8AEs2KvBCK+tXvBSlBH0QbgA7IJ
bnzYFan57w9mxc9kGWUBYeYAh/9uBwP87sQBl+LV0ysYBY7SRc16Cfb4SxkMyEM55Tg3axgbRkS2
21/Nk+1VIaP4zJILV6YauNTfv1S6fZ1JEHbJkVXU0LQgWc/+kW/erAR/IISmS+LzC0Wqp+Q0dXAR
6s8vLUc/4QwX1q6nn9GZwNpBjTV5Jmd3ZJuZt2FIHiYBGuT40u/tJkmA15wB7t0NwmhAesJ993wQ
4rJiEtydJP3vV7fJ2pID1IeRmSgYNXTEyoDAXryRQQPkDEjhCp/EuuJhxJ+xKaYnizG9a5aSiKTK
2PHmMuud9B4ILBIK7pzZfN0bWE1FT5fqs1fChQpXe4IcUpZwdxNsHI1h4/R+OCqEV2DPcCv+f3oR
kcNYUWHLVj70DGO7UhOvqlxZYq+kKUh6P2rY4619eZk/Z0FdLMqEYZ6iOFRpAgaoJ3PB3HiFbbvH
oQLhY5G6e9w17mKxJFtgtvGUCOO7rr/KLo9xls2ZJRW9nAUxtyM9061KACJ4bL9oV2tpRQNGRui4
9/eAQeU0mBlsi/VYjkhDAH3/A8n/YE8IgSex6Tg9/sy6Ay0wIQ3clZbhlGaoEPypw90qgJQyfInR
9hY4O3HTmK7tEJXIDrIzgdngdBBtcV/zbYbrtCGWRXNCDD2jFGEjb5dFEnqkqEPmiFWt50th9Og5
gXqoklxtEr0TMcY4bihxqefIRVlgWlyhB0AzXXLyanJjjT8IlCzoEIkdhsLdKp48zTT2LnpxHfKp
vLzA1xG1Pn1JWzQi/ndmjk2tOiTHNUByz1IdBdsjJgw+zgSsyePoFDEdSUZ1h9ySMpar/ApkSRwA
VGApaYLhfgyI1VBUlGOHqm9Sd51xcuwbsVJQaiKxLe0NcyBEbSuKbDeK7TNU/xPClAqkcGFNxuvk
0BefOjLZemTESteBTzwRH3jXCAbtRBKWBNqWzmSyC3HsxOYSUe1Q4E3lIKmbasHk5ppscJVlspt+
T1G8nGIIdBuAffki8IvXKm+FdznA7j8fbGQT6mgMfy5gOjy4Z/UYwir2mI0NJdLLYkqVicxHKUz5
+1r27e2/DSng8tcSs9eGyQPHVouH7ATxmfxgGrSJFCk5zzTeX2uXFSs4oGWodT/LS33gTZh4315L
9SiUi8n86IrPStpTRKg/1afzCH5VPydoJUyyX2HNSOCR1FqMvoLum+CzfhK8ZIl0MCyfwIdQsxJb
boDCO4GAAO5vvx9uMq60zGChg5tLUtYdA8y5MVq56SVTgBLBN+x6Vh60KvVw/dr+8R/170TrSZ2j
mNM11rY1A/HcdcZeVe5OehF1P4+0iMHgpExqJX2RcAImkzquri5s372tQzlbByXB4f7kM7zX4meA
NiyDEs90WEQUO5v1r2bCbQhemDFfe7l1c1HZNVR3/pjmnViGN0eNdvCfQMonsWWhZA1MLtos9/9S
Mnw+GMuvngYMTPPZy+w4KHiTsHTPU1MM7HikwjfnRuQXkXP3UQIuxxzZoWs0W/EmZiUyazJVy/8T
zG4cm6S2edlqdDwwwDyAZlLApgjMNl8VZDVDNZYb53se6G7+r91e+UmCDs9YUWKM9Epn/otZgH5f
uPk5hduU0jWb2ND3Oy9zRAoPe1rcm7K+icW7yvRbRWAAZX5TvgqPgs86DnaH53PAnGBhCcT3hza1
4Y8KuwSIGQxfYFT+fUvjv31HVHfzOivIXzMl4KDlPuCJE+VeG5sd36fL2nOmzQBZ0eIVxH1O1O97
HCWgAB8sdXbxQ60DH0v3AOUtyn7YgWgBQ1Pbuf/ljl/y9+WG4Z6tS9u5C/C0yvJzOgGGf/gvQsWP
OWU1mN472No3/kZq+utr1B+xqnKnPX422VglrF7Q6P/+yMXaAe2bUMa2IZIdEzf1/jfzoHbSb8Bn
KbQuIN5PU+vqJObhvhyQRxRkhOWipLlcK3MOhvv1E/nXRsCkvUXkqg4M+w2YM3MA8GNGeQVMYJQc
7WBCvaexoX/Sg4ZYbglQShqngzUsFcTypXbQFpLLEuNtAOz9Ha5y0cxF9EO5YpdGUhfLWHCH2pO/
pE2BUTb29P6tWAqrrWEE7dT5d9hrokthe6+N7uMcgOaTe7NBYM5Gv7PN+3BfhZgQsiOg1nYMFwXG
DriSksNKtBt31G2VWLm03tMQ2vyN/6j7DZ8eiMLPdWMR4yOmSH1DP4i9EyskNjrxUhPPo3fZ2CZM
gVZ9NKuX0jsSER8xAZO0oGCx52C2pnK0xkt1rhXar0l4Fpk9g8/Y7yBW6Zuut4xiMLDvXsgqQJwa
v1+NBFM5BQP6P0QNw/NnZHkY+pi15AcFnrhvOeyi8ksh4QLqULIh2hAmVD6aUZCf74W8i0LDeYh5
DiFr/S7FKzRERKg07z2/01AUt8Cxj0rQuXga2L8qS9M6ks35MNPzdBeoypdHlCd69T2kVDqwZYDI
vUg31ghM8RmD1Iuf1yU54sF1+IWEiuljcDhgUDZUwe0Gq3DK8a9LuDvg72UIAxJZuzWmqP2A3M3C
iQ71Z+MRT8ECC5VtNw8asP6pMIGpQV5e6hxjJc4G7AerMECmoSLTaC2xnVgGpx84i3SiMNMHN2RU
Rp4sl5qVci8/JDs0yAAYUUVKM92z3+hHL1ygXZVlqT2Wpn7yPoq1PqHnLnIXetMp1PcouIXPgCNH
F+BFxoCMUDxUkIPAkdy4zvYO6eq1Cg9Qrz8dwKQsplxqIeVbq/hVB8Sw4GTrgJgAXyV94PlTv8zq
26XohemMWuBucm/aTYC5pDl9df+1N9LodIlQcVUUDbZDUqDNuX5opFhE9JistXmunVQojg5908hw
PjBfpkFnsoZR+h3MGdYodGwppbCaqHCA8+XmNtw2phRfK7Sz/m6Kztz7mRul6DP2sVyxRtqm2UQy
Mf4NSqnUlvVWQzKT9i2825DrD1N65/L+9sWBHShoo6JS0xQ8+9QPX+ZNYTR4jEgoRXdRTVmamGiZ
TfeiF+9kVGE03mIe0Hp/OhsdrxTJ2xIGx0TZehOPXD3P9jc2Ju4rhGhwHfF0cO2Ipd6gXtMk4r/6
nxRdRLu0xf8HKlVAksH9qn+KHuoezVlqpQ05fhrpHCg2tN+b6zxBTusvUOuhkowuL9biQEDTsSMF
ysCLjNQ4Jd5gagUOjRJvbSp3s4zGEhwZnTtEXACDJAn6anq06gxLiNXhuvyk49pzkcRUyGEfKfx8
9gH1aKJiKKfsl3ZKSP7sgnvqs6roaOt8h7B4Y3/LAL7gE/8/0fMkzFN6DBnZYsifNb2aCi+/VBTd
qQImX0fF2hKXm6d3er4H1ECUVn4R9uHB2nF1KuNYCAPnG98P4sos7wEtxTd8qXuI3KrXLjdoY2xj
7ZlGIHvwnyhLJEXWDl6L54Zj0dITmuniExoUdodMAf2y6kLSoxwhfoTzH+WgPF98X38VFnwEPT3i
oaHPABlwleeBYsJ+X9CDO/bqK2V7y20RytRn9fSX2sqJ9aqQIHZ3/R7ulOrVtgtHIkeGJlRSV/IV
ISumIDcUv5R6QrWYTbyMxWeNNVVte58YbHPacS4z6DHAgRTxEqyb1+OE3crGG6x/7l0MTIg+s+dc
N8/+75sddgUtJtU86sXY4Xkt4A57XsSvBM8O/yIK6S66F81ccvJ4aMldUIJ7okhKp4VjIUWb7EXc
O6JudyQQjQR8DOp6e8ZV4MG6rcAWNYj5iQ0b4XAKLbuuzBEZmbFVa8KeGMc9mzEQbH9e/XkzePG6
Jh/8CKZUtVDZfj3kxo4U+v8/bpstN3hezOEJL9nWR4/oKD+eQzlk15voqJwLpqZDARLgOlmH74K0
ePeYd4WXl29nJCJKwBSBhgEA4bqEBTTtlAC12PdWbIkaWP3X6sjB4RiowsaANVT8Jq/qDSWmYcQW
D/YG/JsRNUCHTY60ovTrdOs8wn/WQu3tYWEX6jbRJailnVgoNXD7wm2jclpuE71V+MHGwATOgeMb
RG6b8GVgNOEUfNXcPy4auWFtrdHeWhlkT2tdsrCkjRd9xSaYYhWvDegYuSrBP9fceYRvj63u7Nxk
KCVx6vmmFuMoEQHy4nLkEy6DPj55mupIooiBDyILuk3ONkVe9v3+Z6KjgyKQc5p0c0T2JP0Bf/35
FI7RBTwKoCQW6NK1pVLwnTXo259UFLjQwM4GNM22vfwIqUAI2bgMTeEzmg66d2rLWh7No6LkJVXe
rrrGo8+uAbj3BA5x127IWbE2/6Q5qZBPBgGRdWuoomiZEtKibk3qNBfer9rqVkWI/+VSliKM2+xh
p0YIjVKWy6y6nqyK4VvV0YY0NxZ15WO9Td0/vCVZzHCPpLQQVuBCwcYZoHyrEsT8UA4+fiMnye7U
aaRn6bf0Lz0/KHHLyNaOrTLXzwSk4cZT5hVhN3ZpILWEb03Tk56Q4vuHF0AKy5fWsu9/vx6fBI4X
36/0aWG5Otzog+1h4lgInAXuPP9C43FuwQgw6iFGXQRbk5AiYu6/p/r5rH1wuzqVqekPIqOW5hwC
LWgpy0zh9yR1PtvY2JN3sTzsstMq1LSFIsEZQuBb4qj5LzYPQgk2WsZhiIt5eb4B0A3kfL3rrs/1
w21j5EW0j6B6ePUVkAvRvpw0v5eQ0M7IDINJFr98inlkpf2sYKmv77CIaFvCeM3Fh7hqvk8nKQWP
qNfIe0/ut16cmjfjzMvcacBJEqpGe52JSNvtOI9L5r3aud0HI5Fjr7dgMfKcuWDgdLsH5AQLQBYb
MSGyLZ5FZHPe2MXMqJpsO7zW8IuTZZgOz16lFp93HuP88iJWsfvZxYJLbr/LZNthYeyl/gT5HwCw
XRb182QLmfSegkTjTYAvS9He976jL8t/lSHcW7wmB3wvZ1jRMR2uEyvDYXm7XSO4NRnqC/tqxBjW
qsrPrHYR45UaShWFk8+XmSkFw3zftREQiYAQ4LSatBw5zTAde1z2C89RGR7GPZ9zXPxENC2EPMxf
SlHj5apWPfMyBWtVc1PxcZmYwa0QcJIIoefm0c34el+A/Tse3KspQbqsaN0/vgATc0Bn8zmfw0AK
L3l9FI+84xNjjdO6pJfoS8MQ5MakpwXnlGojfYiMQTpyXFM36Jv74NVHEZAmoNVGUIrpzkS/Nerv
8PGg/sVLpD02BAQ9wu0WxelFfkid83aKXDOtx5KDyIPP8W0hpfHr5AFwsHR/3ADOIjItx3THgyth
yFtAUohjROHBnBf8/bbi5O2AOSRTCzra6hukNqAF6HEb2fq+e4rLOfXg5rBBhIoosCspMYHqyv0R
IJm1OZTxyv2fY/caH4ZV3edUsx8FEP27/ZK0m0PtRy8Pqyt4tWqJVqs46EsBmgRkwH8qVXNsJLJM
Ht9cIMKyu0PUCIbouvxnU7dqpY3LaOBgwCdWuub5RXt5B9nI+G1Gf5adqOViwkPdVQwliB+mIU3P
ald8zAOnWcJvo3Esx7+8oIhGg2hJlY3xhe/iKvgzEDAzZca9ZmQu3PV7nIrnMloHuT8R6nTtsHwT
By02oU8t0JRwwBc3VloZ9aEYKfHOQ3PinYlJ9dEIllJ89/pvs1bFcWYTCW831ivYcPKVnawdwEfj
VVOBgCHt6QR6lfYRiui1gADJ5T9bycwdk3tlTNWAcBVxVI30IojZaSEIFf2Nsfn+md3knGfe4J+U
dt7TqazpJvnTJnrg7UAKDLeHa9mLny1iZ3hxefqRzC++R9IrGE3xteypj+MC8gd2ZZ63gIioXH5Z
PfiGYkooecXgP9GulylEZXP5pnDe0QbvStPf1AWJa1Z4PdUxznQBmAfLzLzK7X/6JX954OLEmRBh
A6V2GyzSqhtxmZjcfyEzn54AuT/Ktuz4d/nKEfXP+io4rwpng7xnBPhibPn6cwQccltUWmU/vptI
gBtVgrzGgpdpuO3PS7Oii4HWQw113zjkrX16hYn1vkf741PBebUwIvsifSPiPvB9DTGbNApuLbTC
D6FXzTC8rus1HBFNGeyKQsIswJ/q8S4UV7r2ZKK5SaGgxZhsoJaaHMc/hepZDqu4GfcZfXL4N/6n
uSjKi0XH8PB7eIy7MRoZaHezGNMukrfhHfgbx8La6BPmwsq9v+sHSuL2pJL21QdXBxu8Mnnp0Tpo
HVLjIhOzKiZmhV/kw/0J6Ddpq01R88IiI2kCejIuMJIFOeca1CyAZNPvMwsiviIY9wdtQzNwu+sl
dME8cFWiVT8FvmQ56hKzeC9RYSkSsSqwG7NdjZJhe1wwaOvch9eSGOq3GVhdcsjtSCd4KLlfuXwt
ErY2nlrcHrsDEIqBVcwELF9oKpRbfQsWKcB7ZVr2k6fpqJUFZJFjconmkPRCAgzNdbCRR/NrzOcV
low1rUl32ycUgVNUAItjAm7Pzo/DmsHWw+b2UKXbu+uUPrbpcsGNYslxbGpwRsMhJVrXWqdMokXL
U6gNO3f1KUI+3xuNLCN5Fl/tkuwzOCvYdvJ7D70+mMag+2yzAGkdG3BnK4II04TwXqs5eTuSzplA
6VRAZ+MN6bsk5TPrYYFLw+BXMkPWRPrGVkeS2liAzftwEzEg6l5eAxJOtxO9MjSP9y9EPK8XMQr8
IjB6OcKvWpX8eds4V5YxwIl8MGIRqxr3TdIvkzPGQ2p0ZUg9yuPnzkEI3jvWm3pgCbkm8HYU9sFa
VdtRrCMMeGafzENPoNi5PuyKg32Mq8jwnyIWeDEWgYpq7xKBIML+BWK+9lNE7FH2ZcHNca472e3Q
dogmGgQF6+wOGvbIhPlxyVFVrR56G8TCcnOGK7kOE/PrnYjE+xJST9Q7iN/V7PbgcPdd1c+q126h
VJDgW+PX/uNbrs4V3UlaoopmcLL/Y1WBQndri7Q5q+LZZzvWv8mJTex0CyyA6L2cBcBZpwz+kLnh
H1p9/GysXioytC6glR8OnQG17kG8fMwtdJloRnuCRYCMRnC0LHuUs4Udx2tGxM5dZ7FV5iZ2E6bM
9EAt8nebUz5G8G3Iab7oiLI7/wrHx6kX+TZxnHEiooUZaMXWrOj4EJU+7O6ekD0hOgadMK1j4X28
YSxqtjKweeoXBZ5s9+c4ZJTU9GVhVgn0NtKwinm2Y3VVPP3UKVybh4lL1j44/xDUCDwVzFm7gjeA
6AB3M1h9k77RSLsQy6PMU1QNqHVkyKTMTMu3etJM/aLa37jx1ZYLR2a4c7+UKBx7AFC9NvV57CW7
rPXSJMhYGOdAeqcDb9da6BNT2R6Oe/4wy/s/ssK1OYypn9KhrfpSLVhGVX8WsVu1Aaa2pihny/El
J4KCudgSSxozKgSzy9aY7bwL66Bu8oIlrlXavdHX/myc6T0BwDm3t1f/kawvBrGSRlw5lvRJj6r/
kxC1Jcvsz2KclIn1Vz6+EYsBzXmfpQBLjbo/fuZZDUEmG9x9c6eHtT1n+TNHMBF1eZwurDNYSZ5+
TgKx5huLXolapeiipztanDihynScxDt8n+iG9x5jCf7USI+8DaXyZ2rWwjZ3UDkK9A/prDJiPgY5
dH+J7sMEO2fkxYC5Ascydj4vcDkZbtPwWhhsoY7dKqv/DNu9/iufVpWZXnBhF9sLmcqjWqcRyFJH
TCBQsVWJrp//7Hnd9Q51lXjAvZ0rA5Wl5YszWjGhQYrFvgEZMZrxJneAVQAIGZaRNhef8UtlZTZ6
KmW315rpmmkXe9cfcPzFcuqvXBcUkfi1GdElRsEHDSXqY09I7c83PLnavSdOnZ0xhZFPlFND4jEn
SUVp3sQw4Un7ZB6O7YmR3zz9i8hg5co49rt79GPWBGupXqXzgOng769u12DaoD7NwkK13VsF7EDV
n0Ni3xVR2IyHcjynyDoMcOl3ws/VCyOVxKjsSANIFc9BnsIZgDL6nYNr/bQ+I40C5qWPCZLnznGh
whRdQeudzdQgV9oJnQ5Lnl/JfRZ8x2JmMaVbMBK1q/gJN9i8AH6rEUeDSTUfNPmuN+qKCUy3MayZ
yTtZ6oERSjLP4gILlQAKhYurJKYLA+ZkFej8jwi6n2WqEigT4OdzF616soprcxEYTcdndZiqU5fi
cXrzptvqVSGAAxE1vNZ71kcQvPf4gOEgA+rplsDaV2ZmOxrnwkIQ0NG8jH2A9SM/UCGQon8/n8xZ
Cw3wX1F042/8UFtuw9QtoYXEe4b7viPDwjQcaqQHMV2fxAqfnru2+OMM3EqC//E/KDBB3Fee1Xsq
z6GS5bUzNnBx8bFBFCm12HJ8QB+p/ivUoAdMzleZakBs8u9QaBcHCNNmJbXjY5qzNT5Qaz8WInIk
TfEs2DfjR/lN0t2zMGd5ElnvkpvBKLKAL0ELjEid7nic8J4ZOznjsF6Xmk3E5mylsh20q2t7r8EC
BaJCmmPcJzdf3PCD9axYkzBBJVARqKK0kI+CaZ2U50yzdjfgYsfDMQ4T/YkjgsTcfFb85c8mJ7My
+MQvMH5nD1m3Vv9FcbroVuQbrH0Biqhz6zKFax383wkpDtEVUYIsCDnCRxMcHk2zPtdLjkrBo90/
q+otTFJbOym5FDOo72Nslu2EGCWwWN6pGRAqil8l7El6nictaNrZu6cfDPBGxAMnnIFekVCNxxmT
CLYnnxqR1UL4cc4oRnnmoDkfC6Ipd3uF0nPIKfcKHWNgrycJB3FoQCgZYRwg3BJf+KdZavPqGKOt
0//w7LQcYZKnVKgXttCCJuvoQWbeDSwIUyV3AOtGy6hwUIDjGXTOfN9AdSZD8Trr3wwC1XVx1oC6
y/qQjwaEZdNUBG9tcnGqdr/s3bCDjkrl38OjB4QbXiGIHYlJhokPreRtyO2S3Eh0qfEQEvTU62gv
+PBU47C9cEvkglhXsGzJ+zx+2dIarMvfFczhmDrwv4d3ikWxAixkYKfwXSm7MKC/UxAV0tZ6tBlN
7T1MUapPe94OHLLzJCPmBhHdHpX1EeByKy/z5fr8zvypyOUnjEo27e8bDQbl5g4Zb2c8WJ9hBsGj
W9gyXgOUFdywae1cNdzbnplwq3wqDsB9LZ/Qjn+kULhkiWD6XHwMfPIN4CbkNdMFNXZt++YQmukf
ezYo7XpWHxxLIEwWnznr8HJdIbVblSGdjYGtwZZOu2p0lqkcEJarvg1hUb3xilNVICwQKlbu1DSm
M+5bIOts117A0wbVShQ/MyTob2S6YaJlMDyBOIvhSmqPU9+G2ZFRt4Pix97E5tNvcOQnTm7zDBVg
ydRUwzT/Wu7aSK9afXT/VXacAp19Dvge08BvpRVpUs9O5ElUatkf5CzeVJbQJsTyE+jJPNBkr4M+
U4oO+ikhaOCH2VSjcsJ/HUKnmtMJRgICXAhEWaK8aREo2E6jKcDvD2RfRLMSF7CF4h69Nhi7Tz63
wucZm1akCB6D4yAsCfsSR1cuPMF0lWXLXvMbIFAJ7T8iugg8Pion6pcGTrBLTiEry1qdrRYNN1N3
m7d/k3OSGD8QWKN3UaRI8zpD44xMHcS+1MU8Wjyo70slFZQambSEdwCQt4mqWI6XndeoV74mkGIU
iF9dUbq5UOuGzO+c03I7jMSjSU2bPtWKo+wxFNCoVq41AJdJM6G55vCqLS8TqpDp3HphvE+JYP1c
Hw9SWGIEA+aA/m+lt0IF7t+OU/71XCs6ZsCiFCDaVFHspiapAgYiV1P7MwU0MGJKSd/7HaABopoR
zGN6madIkEP9CYCPB6tRIy/y55uzkKOKqWTM+KMbI+z4EeuDSGGc+3ffEinFlzOPgPpCcboyq4wT
RxxKTONkuV+IcvDEIiVNIA6cvjP1lzWnyFN6BXHK9bselYfwwi4sQ5RNDJK9IFCzSpOPIrXMIS7h
i0sGhPXol/FoBSH/nmALDeu+nD0g2p0929NyyAZE3ICeK6KUoX0Ngdu3De6Wvj55d09FN7VzVDcr
VZIfInEXzvwLSsRKxMMPYr358P0R0hlywsrTSKRwXVC1X6o0ruPxcARtInVytkz0mfhEVk/ZJ2ZB
xFePsy+wln2nu++20hYAqVRdSJLKc+r+C9ZBe/djXajapgKg5ehCVBI5BAD5cyHxJVZDGmVRLQaQ
BcFhMe9CWvs88g3ld3rPK28WpRznrByoxY1EX0sNLV/9EcPiefExyRGuBInOh5FhQ93AU9/NGc1h
/xcXgo07Okjl9OThzFLkVhz6cX4dsYqdXrhnK+BOxQgxqYTTrL9bBCe+rusOx4iy3s26U+0y63nr
sbkPM4N75L4pHBKueYIJ6gniOOzdyh4rbOunNLPZvSIj1DRqkq5QduQeAEJ/9QXDEywZIL45wl1I
omMyh1fJJG5SWyOyJZ/DEb/IeZRXQAHVxCwNE2siKqqOvVP9VHnQcgbxK5AFtmZs8uR5U/Gh9UsM
OcsVK0tf7sJUKgLJ6/coITpYAHjLBS2Z7/91CVxXAazhK6Lu3tEutG7nnW5mI1oW1MgSmurjXqpf
N4p7OzhAblSYMSuiHkHhU18jUYHgT0m+2VWptjf9izel8GCvB4qr/7Xk+GTp3iQ9hahBftPPFq11
N/sNnNLGXOiDNQ5SD5UAYOwKmoKZg8U0ASF3c1gcV3Tox/CLqSI0v/+NYkSdnXVLIxRBekHiPyS1
efYfHBpuheAItAmz84na0Sp4A/c0Dm/5GUSr8lapGa5OVdpVWCZ7xJsaCBgLlVHu6DZIlAMyxEIp
v4Yqu5KC3z4I4kpMjiXS3jc6OPgAQgFKTAANH8V81PBXIGwQFBRA+qC/TBhn5E+w2gv5Eyg5TEez
z1RHJfEZBi7nljSw8aWtjV8m0OxEMcmRgHzUWFVUvadFGYcs7JMARhpOzvntXHxryrWtzQzQH8qW
pew0hutn0w7Gvxv0ETmPMEPzUM8/msvVQblUpfn+YLhYprg8Vqy2hCfi82yb1L5eZXeJX1ZghgZC
z+QB0FlXQ/RsTgZ3FgD3YmuDrr2HrG5C8s5+P9dfrZZ5XMLoQbxcqCZudHNIVf2jZ4JymAZPS1hO
IQ+gd3oqsrxwIe8ozhajc1XWMqnXjqrVshUej2ofZSDT+dIjHY+TZVKfy3aV/LDP8Z87dHks/t6w
P9Le28H+BTrsSPRVMeqWQ31GahGs//eMg7AStUYfxE/nOgiiofLZzGk3CYI/x6td3/yPQf6998Ob
M+ygrgiWvk0OINIpl8MONptJWsUAfEeJ4fCzC1/wgHrAXsOJwVQijnKDOkinjgDSN1Xuj2ZJeVlU
nM5d8Ni/7ilxsP6w3WYwVbdrzTPEY4VNr7Ed4A/bTGDGmNSG9Y9vTIN6uxuPryZu4pZj3vX2HlOT
SgfTwJAYQelg7PezkItB1wO9lJc1l0QlovNgLLogVW2eICYjUFm6dD+pLx9oRB57jxueXXU9rG/a
RjpklQA2fJcVO1jfE6vwWH309QlQm/+8wwK5T/AO8N3gE6jVZGSEaPUm5XwQFgmnOpvC2zM/rZyO
TOOzh/0/UQf1H65GIpiQuTazt6zxm6FYcfu77qZpkPK+8uQg6XILc5gzKypya0afpmgAWji55IcA
Vvd4NrftGxEWGXoYdMWlfj3pNKvbLIsSmHsJdwEfaEnG1ZrnEsl6fgq/k2w5titf3g+uTa+5ZWxM
+APZcJfz6VJSz+Dkaj58ZgdmM8mYhmE5VIdsOczN+iZjyyEVvI/lOceJG+QCcToQy1mTmPpA3E63
KIQriCaMTkz7Lzvg99hYTb05ckkCexBEnUeVfdH71ua7f3tXikrYK35dLz1rPnqrhLqJwQhXB2Qh
YSOnqu6FEXAhg/uQ3V2RwMTpPdepYHWvhkIf1iyzNPhVI7EytbjETpDj4mlps567pnBIx7bfvJiO
47Qzt1ne97o8/lt/KsEzuiBpQGmNQ8CT8ZxWoKhPDVDqNpnsEgOzJM5tqmcKnkmFtWdNZhvbByAG
vD0KzNo06vGd5Bx6S4xyv8VcekFu3BtLrext7Q+qfulrp1vYsFsjFAa/99o0JCO+pYArtvPYlfTe
ZFguJ0vKttYLTVC/i732NRJXXvRLcWLH/Bh+4refSPlLRdqa0Pfv+niO+NFzoVdiqnwe8/x1pVpi
ok5xVlfMPzv7kE9KbdJxxk9WP4fvX/mJ9KJQj/p+qKA6xHzTPvYgGfFnpVufejmddch8GJi9xDzx
T1jhFPbhkj0yQMtA5fJKX5cLR7o9qZxgRx5dPDZEdQhU+/lZMxtyO3wRSKLo6epNMu1/3bLlBioc
DaBGG3VocflQs1Y4mhCwQ8fJWe4ZSfkc35Gy2xKDCZ8Sb3yLgRPWOfwTfyDCncJDoDyaPEr7uLWq
ZokshTCIaIShm448674FRoYsQyci7sWijUYoix7xJem1DZmImf+TxATa5O/hWFTyuMhoCPxjUrW6
81arFF7gUYfswfprZiqGuy8Kh7TtxAP7CewiRS9/uhKPWVTRl6eYpopYxhiOHB9n4HgNs39Mix5c
tQMKrch4caojpE2qO8D1SKuABeHKoqlZqIavAQfLYzpFb7XOz5mfkJpu0Idq/9rSrsRCScaW9n6B
3s7VVMMoKHn9738Kme03OKa/CsGgvitgGMYzqUWT+QM6LZTdkm2wMeusDzFLaMfArnn0m/fhD3k3
EDMypAtq/LGyeiRs46V+WgxR1aW8WI1QXoRd5BxcZkRpenwB0EFYBqnM3FRQPFHDTviyXC09Wone
RDY0IMa1wEAeALehPJhZxF/IAN7CcpXvfHmRAsT8VmTdRE32Lfwr59qaMPSg8UK/M0FulstTni3Y
TFqYOlz9GXcf1OY5vZr2kREAza6sB+4+4MMQ69WMcIZLY6keHp+q0eiegMLkvSAhzHbjG0cgnTdn
vADF0ETkJCv6GxETAy5hXacJ7i2GWGUPPnJCfdU5UDWFEuZo+CF+2QcrQjCJ/NEjFHD9eWCUesuW
EXZ9gckUZaZNSYwhtu4l82WMOo2MbSCm0SNlIT40UjDnmaxJ+K/p4g2iAkx76Ogy/JMk58D1zlho
gQCxOXMlb8FV1EGa6MHRYansu+8KRqZj3NMWL4CqCE+g01nGHN1m5D8+/nIAn7WmdFj45U95nLu8
vJVqi/LBYXOplgZ4BrLISw40RryxKqn7MsympakWnnZnxyfENBkCVLUgLDABkqzeJ88DMuNT6LF1
xZzjWcwJv7yo/rKTGhxITp9jd8iTI5sXXxL7DjXaU3bl3r1lm8WDWZGTqEzYuKWG31PYXGTiya99
TrJ0TtS2q9yVma0gcPW9E129+E5Y0/+ggvDXb6UTnt1Ph77qGbQqFQLKdBSSXSxBOBmSCqNSByWs
2ezqWWRc042rrFwahnC+TlSTzkwi30yV/v1yTeGza8jMTcs8CmPBURb+kjmpRg9+Fi+WL3lokMax
wcXe5R4Re9sfXO+ciW5x2cqU6EjHfep4Zos7ST9AUhIoL7ulb4R+VawtSSwkWv/Q5chbvE8hRLar
RTrS1XDY2lRhgBArioOz9OXGKHN+efPERptbhN37+HP+eyxqpI2B0Q9Pbj1azTcKgDZfH+p2ivQQ
eaE0PuzDmd9RIgyNil0G+agfZMxy+iSwz7pVdnfq/YBDdmjpC7HgHrrSCy8y3+QsUOP1JEjSPtIE
+WH8KxE+b8zKLVe0k0J0KvF2ol13doJaoJfPo1qYXHqay9owTMls0lV7kv2suLyDVgx23m+BdHby
UHgRvVsYwRcLRcJPQI0i/Iq9Xl4mpEzyacqh6ishBkjYmxJG5jnD34vnvDoel5w5eedjaus9G4na
9XRO6EW90SW+4hsQqTeGy4/XT/FN/7+7C9nI5gTFYI0i+7ofaRCXTFV1iVdI2TkPLOi3cn2YhIY2
Np0R+hvPtImWCdZsx5ClvpBOw/7uDPfDBhmxXfQEttSgexDE/FkSnDDTIh55I0xCOHS5sKAHFQL9
glpgFPmGZfzP850S4MmWMMcs9ycX8NJ65giaa7cYfOP767kVlE6EGHR+t1Tw2tqaDMR++lPV+zgr
tPF0savmEOl2hgOBc7YpI5LihlEhbCXtvzb+paiqw+ei+G5p5Tbj4ysAs50zyQusKOumEKG7ejGd
gShWoLZFqgj+O2z19e0dzg6X0FFngYjwahKuWVnh+tp/RKuu/BGvcilN+t2F9IKwCTq3svRtSIh7
+Yf6PhxnAkERy8povmPMFTZXO7MHdMx2r6pRzPoaWPvX2u9GhVwVukMAeqQl5ph1nvMAVwXmIfc5
3/xRYq/fE8cLBnsbonGd61aL4Vz627g5ib+fvl2sScvb7Y91HEW1guoVtYmn1oDJ2H4d1oykw/Ij
wv0vekcFtny4th7ms4f19lxl1+8hZ19VykQPuI8EM7yh2J09IEfuUi/ZI5JsPJrjCZ6nvU7nJyag
fjcf+2WalIqnAyO8ntP4ftPyg9AzEmPVK41QnZcypW55nflNBUdXZ4THUGqjX/71inJndD7FDMZA
JJCq/xtfHJTRo4mrHjcV2kZNyaUsjHFOWFlzgbAyUV+slSj+Yciv57B+GPST0dQMVOK/gKlU/5XO
kcfIqyQ9ynLFDZ2YGeJ3FabRK7u1xl6BZCnwHzPtxZpQxCdRDrtA42M3cw/ZP4siamwLhsjYXBa0
AXcL8lgM5s9JKP2+TVwHGFGNq2x5Os2njwkMT1j28A4ro6UECylZKbz0x6t3nGWFFJq0XehrtJeQ
Ka2kaiP8aevItaHIavoDeh/fJc5NImglbI4qLnyhZe75Zivp1yWxZ+l5AJwogx94tWr6+XTatFw/
UAmWnykRj4FetJWwXWVbzSxfz5IBavmmkHD6e8hUwcntxmlf/wu7Ocn0o3RttX3mnoVeNnGd1C9U
K3vdKExrRvdpEMu9wAO1i3eju59ZfnZxXYOHywsKInTicjnhpHZy6lpGm/QhFIR48FvkCGJTjKOd
zkIzrJaTV/lchFhxk2yY2318h2p5m3Ze6RIkL+9l1mpM8koUzEpNVrzrvQSmF4cbi8KpQGYrZimo
WGZYWAESEJnGSnUloKepuOlty48B7ArmWU9U5asDS5SFkyk5A0fBjtXS2L0yuaiO6yFzSPpu5S+v
dlFZ9SHKlxVXTzKpQk7UcCjYIl+XZ7CvlAU4lP6fvfrzWeUhk8FwQb3o5i24vhcfm23gduP9PXJ2
G95HOo3+h1xFo3uaPouBQP+vyE7/uy8kYrKwy2YN0pCzRGvvpxpFm8i6nkL2GxGbjk6aaBvQw1aW
LczYyuYkoz29JGzZtLk6mI4Eq7Kw8sU+2zFErio5GOiaiUQThrZd75hn1H/cRLxsC3An3ZDqdF2u
ZpfAJrSlq3rm0gkC7Ivw4Ctl9xA9CtP+nN5PMvAOXkVR+X2DfsnMD3l+6kmY2gQNP4qd65G2tUt9
GjrviFtDd5EjcguvL77UnekQdvmEv/CNaFYhKV7oZk+so2nzYLhMN3baICNbPHXSFPnZsyAd7cEN
rOM+kqNo5TtF6YNPLVb9Cmt4PAjRD5xEprR3QCXYW17Ppl2sGPkqCxUargmH/erbKz2lsKr66IJf
SdAB1r/j16JF8r+9h0e/EA4549w7d7KirYSrrNTTy4lbfUWfkf0BjEsSY2ZJCFlwgkTV2bLEkpFu
gDQRIU7iJ3lXeXFOb6oRzt0kn+fME0jMLDitREoJBM4w7UY7fiWLyHuYKQlUzlhh6OLhknTIqNJE
vp3RjETgU/TGTzy0AkdEmZABUMi5yiBGBbgvbkMQz6TM9uXsesoLvIRtU4DknPKC489q12jffkLF
A0TpRWI/WNUgywwG++ZhJ0alPXPKtfSfCGPu/1oUOteg69E7F0t+N7b4vbucH4oyOwDmBF0Zo6//
kebk30Pv6VIm5xktwYaumQnXk39ZzqsK5zRQ37P+pQ8MOG6rGYcGLwtgCZEakkOU5eyvHNE2ZJXX
XdfG7cETgZMAtUx9Y5tQ/MHFrP1JzmZIcPI7PgbXKRgqgQMhYdDZo9pIHxfJUYq2qAAPQLkBqjW4
GPc867PH75XuEKvP3kupQSVGhA80h7bWmPdrHL6ElFG9Pyr6MPs1Gzslsm2PN+LWQlTmld2vtJPU
iGmFI1EIBy2ank16eYVz3y63VRK+K3yDRrRJeJOzpm0a/fBd+VmiULFGthIoBAHOR3quRAiYHXlJ
7hGYX1RLxUO7AIPam4EvnVFzgQ41gbGXxpMHZF+Jr8+nTr7/OrNbWtd8sUGPJC4EgmRyRr1aC03T
G2ffaV1Lt7dThq1CqcCrHNqxOaNEK1GVWOtJc5jENF/mmHNlQFT2TUCgsURl8f2A3ymUuiPiolDq
iljVmcqO+Z3TWzIFktuWK21+gqWrd7KjiTF0j0tWe+N6liu9LGJQVsRehRvyLAzWcDaOG9QHzmBK
2U37QOEq3tfwCsltHY7/3Xv4RDpWQzi3dc4rr1abwqTRJqTrM3BbnCPh+9ynQg1BIRQyCr/Yjvzm
fsoEWVpAk2gJqZFC/NgupDrkjuATNpTDVTgW1t74v6EMC6tf7u3AS5LuT7wVpxSST665rN941mUf
migtF7qb1uSeyRMfbvtphlNRHdTC8CqxqzQ903ASkFpUhaiCnKkbenZdPzme3aY9H+4E5yETOCI1
i3G87zoIg7SwNu/dtaEHPB0kyqfpNZCVbyTD9wwIUKhxGd3IKJes2GB0N/W+bjB6mYfsQHQ7VUT1
8jBnC5KtWh29jgWw2ajXLMqBnmQIa42TPXtPpGZSix1DmA+Fl2N7efEJ0Xq0yeXGiKG1ek3tegEF
FIqHlRWWyoTTFlCAJJkEc3zvf9roClDr8N3NPT50m3zIA5PakVMMhOUFnODg6FJGhgmrfsn/BCz5
f8EO0Z9KT19n8sClJhbRRFQUbMcRexdsjstp9J2u5HsvcMGuYcq1J4lwRrn3CMPIgUbq+Ze+GiVv
fSN2As5ZOY8NzLM/dtkKjOwcN84rEHCJbyVM3cr7ay6LvVPMgS/5P5ozXFN8oIxpp3PCiCttEKgE
OJdMS0TbuI9UOyYb72U9mbgjx1DxNM4UFkif+nHizoyorCHlavIM3/JkJas5co202GSS2X3sw9oA
eh6mfcJhbkidfk+k+xIojsCvDXpfATVz5WmzowKyeWu77mxs8ZPTRe2gekWoxTAF7W2logi/aNjP
g1uz2pJEGLYqzDUdw45YzEstoNQiyg5CFANKuu25Bjd9OTAHE3Vh4iVNQbm1G0agNG1iISl8ft5+
daDFrCI+FOGkwfghWJfggl86obqC8dEpkyUhSMSye35Vv/QMhrRIqe4kkyG5aBNYGwudRFimogy0
1F0PltzIIbh0tuGvoOUjh+3i2Sz0F7gmWJk3h9zropa5Nig5/zwJfFXviqkpeX96djtDAtii6YZr
GDZReiWYlcZ/pHqIbyqVddpNV2b8eP2zW7+jnh48newP9/iqyiz0+vhi7rNIXTyUsHN/SGLMdpgD
bl4DAjcnV393ySzVh/5ikFyjro5YhjUqJISRC7zk75UqXu1kOYMPC7mfJ1Dy+LDPPWPxqEjQAo/Z
EXntpkAGW5ywcMmxIXLW1MLKIfiIZUCvLo8LE2fqLNxN7hxneG9Ctq71kZ2moWXs192xtUuKnH6U
y0RZKe2Z1LWScL0pjY0L7j6WgUnz4DsKX95ZhgI8OlHw01N5jzVdTP83jVTyde0iiFXfLuorrdXL
3jAlmDpWVzlycdSyqv9D4zTX/xC1WH59Pl6tIY54VWgvuNGF7qa4MYDKZXSwp3/0g2b+xVFgQc31
vuBDkSyMimDXmYYIM62RQyIokW8KXo7V2ksqWMluMadv5HQv6qexae3PZLwFNQCNjfhdnBDeCyKl
Lo2v6Fl8I2AINHqXhrlUHdF0vAK4EcCDFU1XMLjR+w/RKDyG4vIds2D29n1ysukMRgGuSjet86CC
PW9uAj8KdnQYtk5TMr8vbVlZeP5L7oyqNaTpm5b9UDs57ly16z3/AOhOM60F9bSWo5dw38TyJcIJ
TZNFQLdsFz/Y5MjXt9w1pu0bK97a3Nk+mrodXOKrhA8cO29eqw5V19QcwedleOrWAtOfMdYvO+Lr
a4H2v1izZglmk4NIYBYLlUflF6E0RR34avIlKpvbVhfBDaYvgUeOLk2cIsKsv/Cqve+jQD6towZD
lldeC1PRdoNrarUZdB7Q7JaBxUM5ERtu4mvJzmCpR1SCYsKK7pcUw7JiCz1PxQXlB9IXz/M62gZG
mGF3dwwtFjUs8+6DnQygAcGHBQMJJFeXMaaAhhgaSr+t53yhFm60I50RxzfstI1Ro3SC1lMUojA8
a2RC68awILaCQYXaJlwPXjoEAzO5M5vDArNr6Hsg+qnI9M+pZwAWDRim0rzdInvkIsRy9gmHxdJ8
zspwhSE3TJm2Mr9AF+NRqk9EYBAd9fOYTayRWDYIl/NSv9pXHEHbBHkDlcfcM9Q5Fcq4RvRrMybP
A7kieygqwg4hOByoywclgSG7CHXVxVdslpvm3nUvloLbBU6Yior/a4OfWYxS36+c0bXgLYHILbdq
a/xrJG8zaiYI7csSqW8Df8jIJ9pFLmY0ZXAviij4mUpAvu58Kv1HjFRXX8G6NNBpvMHFY5of/quk
LxsutG++MQd/FjvpfD9LPaJ4L3109WtaFpj4WwQaN1mmb6aCbVuWNRzwfI9pvVsKo26NtJIPBkNI
tgia5Rx23zNC9bS2dSorue5TQf6R62CTXaAxthsgMEbFlUgEbTkQPnFN3jgYPn93200879XuUBoZ
w3hcG85al5gk1AvpcO8oMmdiv4myVB7yHsXFrjuLdNW7nxom+C4i3jBG18QEqRk1L13mBzhEB+m4
duk6IvD/mO6XTACaZd6XsY+1Ftmia/6XfduPrq+LUOhJ+5DgsPmejb/gEDCS57BWK7MBmyH2dwzk
bGOvhFztAhCeVoSnnuBevgN3L84N7RjVsu7zEACYkoHToof37PDXVJlho21j0o9VVfaKbRZOWJBe
U53UgLUfXuG6M2CGpbqgL2GFJBZiFv3R+FJL7q172FogsZYejvYwj4gxAVxZfEHlzwuaaqbmBwu5
vfO+jqVmTiMI5PJRiMTbk25yI92RBRTeKb53zjfLlKC0zSE5VBSPm8dwdaSyIQpgB7YijNgaLFJA
8mHGpS00elCRRGms/jBCu3HASoBDsmRpDhetq5vw8GYr+7tqpwIUNqI/k4QRDVHepUxKLOZl8c7Y
t5XBmPKJxnpneIwo4FciSfMxcyKZjApRuXieyFmtxdiU+IGLZrCQtdLSa5aT4ix26jybZhoAWsrk
be1YBSxmXPBXKC9wzSnFMn7DnvOn/5ePVE+N1b63wGOceFJDM/XYChfm3M6qiyjYMGMUHK2flrli
S+1XU+8F06/MiOs3NOo9MLeqOkU0QWWMNB+jF6gUfziTDwqcQiO1QzGfUy43KxhAd5pB8Y9Vwd2S
kj2USKH2EctvvgN+EBG/e48xOifoJyVFLOQqtTc/h/cb4NU5L/J+ls3pxzA/AdZq2/Rl4dx+m73S
kJY3rdRtqBGUb7v3XbzYghOYR7oCfmwvQM6Q7y+gPBGbgkhp1kdMVK8/H3E9R6dG1F5fgEVOGmsy
rU9AY0i0GneqkKQCx3qK+YZIWN1BmcORgKkiG5ZIKbM54Y9ZDZpmJR3GYRVYwdIHT6xLx73IFowv
aIRJxxG2vxm1INAWY4xg8PDvdMeOtChbqkiYctvciuqgVhu8F1fkbi73PMdYmmfalouah2gvNHwc
vbu9m7BQ1HbmUkFGs8HpLOQKmn4S+zP6x03BwlmMTg9ixMnbRbO5FYLNnwmdybFt6Bx13EnWCltm
xY7V1qUEAfCI1x/KJ4x0N7ODWNELnuu8Fki8Hi/LB8VZGS7a9e5/ih/S4ULjDt791r9shiYaQ3oG
KmU6szkgGyrC7NMCySdeXVUpqS4gFT2TiPcz5Jg2dPIxHPkGnzlB5ZJqWOU5+X+47/IBS0rpAVRB
S2WYfV9GFyBC+RlyKWzIyfCqmC9J300J3dWConR4aAaa2dS6bHPfLITSgkVleMmde7fQNzw6r020
pry20K3BXREEK6dF0+fzaz7A90Ed0p1o24ii2+AYrvaMGneZYKU04v6FSlYbJ/T+KvKn+krv7FSt
RmV7PAyyh8g+tLSvr+ohw0TDoJloKPV2TpzSpyU2plbSIEX2xBGcppqC5+7JQkxsu0F7fECLIOmX
qLsW3CxJSP7pBjObvI21v803klTlXVCooFOafrY/Xa6TuAa9PWc301QhFFD2u4AFISelg4vfW+Vy
Zu0xU+LWOgC9XRvjlP5+fPMB51Tim9pAAuK9U1JmdDIGLzBHYYzOHTkMim+wM350gOe07/6eKrLT
bmQEq35P+XvGuA1/Y/ae/l6upDow5p4xNigea8m5s4WgwJC4I7b0xEq64TT05o/cgZZ/g4zQ7KTo
mDDPUvVnjjyntmDRLbnTyNuVKuK1q9+9FsGqPxutaGGMZdzcsD2O5JSDmdiF+iywUV4b0L5u6hff
62fQ2YQlUrNyswKFmS+YlhcoKb4ljnqBPEZSOve9EBRwbXw+4hMPaVqdAzQLS4UrTFidOX7hOKQG
izAUeWPdkI+M08pa3vlWxDuDks4S+IHB4J3Y0Rs8KJyogRHvnKHm5uMfXG4fA0WiDQhfJykQrACJ
eUS3Epxi8KNa8NIf8h6OLid+KyNIyDlqXdeSdrvy7S2jNhqpLNaFANds8Dr5RyMkvFKYTFdI1Yem
ISskqRIo1f/tGEJMhg4h5Bb6wisW4JZQyLlEq8zj/n1PfLFWXXuw1yjldqv/OsQiYkY/1hTnM1V2
JRCtlE995jNeO6nFNaw/4HBBu2CEL04Dhak5PHzpkR2tapliDVn8J4XhXH8Cxel8ygknexoQNK55
YTDIJzaD7VWOChD+CZRa5qPZf6fFOjotXgucHEKS4KnRAPPbk5/Go1Td+SRsp1l9aoqJqq1xClU0
KeCAo6xJVISCIeQZDFxTMDFIvpepHao/yKBWI7IG8M3Wvm7RsC3YP6e+DvajMA14kyowtwQNslIz
LAIfIeHIyVMDxbKq1tTpsY+GE99qA9zoi3hKrLDPsENQRltk8+bND6UKocx+xELQZsZDWWtWTGrK
ejxU0nwN9UneUag3CgbzKBCnxkXOYnEIZL5YQgBRo79l/qIkUuazvo6aXMnFDsqPqOm1TZFEPhPD
4NJ3zh+Q42RyrCEv7BTf8bvm+VwK7kTK3uDSBOyY2+ckP4In73TZxoEDMwnV8N0jlPHmwyMkhvMi
csHuPT5vfQ9/zBrw/A9xiTcWDpBdw1VOyJMfCY2H8jUCPgRnL1sN0N4rDYmoGoybhWzK2cznk9ag
vHD2Sbma8fLrZJ3UiesVgg52jlxZld66OPv/j0NeZApWtYWFKaM6bf3h767LF0iQpnp116dLo3k/
5McjOXieQMTdKqWKYDMvOpgUXmPxIMCwkhzBbUJ6r/es9XO86W1M6UNa08lJWZpTzhKG0AwepFls
CTvC+nCGkWso54PmmlnVtpuV+HUIske2iy84cntgc2EtM+iyjdnn6zRO/a+SupiEENviQ5yAEMql
jju+Xh0t/jk5RxzQ3vz+d3t/eoxTvfxQV+70ksBKhsE4W95aM0Go1xUaz7ELfNDCew18W2DXu5Nj
BAIy8oETfD2pV+KxQkGJII1PunJQ7SVNnX94YLZfuMiam+OfX6QCU5AKa6vUaculKU9BelYLJWDi
VeIs5cgSmpYFat5KRclOm0W+ffab1noayN8DPQGQi9LIWDpW5wXa33rp2da0qo9WZJhSYMvCqtKH
xJDAI8CAPYLz5VmcgdWns9IWHdGXWi+dC3Er7olpM9OROVPutiCMxQm7Anhy8N4ExxaMIdItSv3d
as5Px4KUvTAV7mwYZDJfejYhf0q6KTvibG/BXzh2NMq344YVj7dz194mMfcEBTIf5P3hkuirNalT
l/MG/U/9ZAF9weMV3X+p8tBorVlEos7bCMwDDRQPQIjfcpgjpm8DcOuNVMVNAfLLpCkw27nqmQdX
56yvZvps8BdnPzCHaGXALu6dvU19qLkTiWJaMaIrX8+/qjgYQWQvck0j9uNgzmhrwAtHjxveGlQQ
N+6YI6RT8LMjW2UHXKoiiEgAC5KxYMZWOhqhGNBbkExwcn7dAqe1hTQ48IftlG0IO2BxS/jfIUZM
pcojhLn+rp7WJOWpwHJUOwJnFIZuPzprXyHcW2uc5JabeYYpiIZwEbBP9owVBp39KJuRfy7CHaHN
Mw1YP+a8pDoyV6cVrKWXgs2WG2UYT9iQC/vwOzubErsi7zPIMmFDyPq0Qk6ClWSfpI3zuoNeQ+pU
21m4ElMArilIOh0KGKbBWL2hmZLj6YPeZ2HO0UL/jPUqHx5RluEiQJprYhUYO0SZDGcZnAbDfiiA
Zjo6j8+Zx6NvnLR8GmU93e/ZROnd3YjUDsK7q0iDcZIKZvVIHY2gsfmCw+GcyvJn1sF91V99cQJN
z0u1NaET4XxiaE9RoQYzdgUp5PrlY+iQnVJYbhQ4zL66cXpqNC0p6fm5pg022pFBk9bCVzlWY5Fx
ZlidJYus8hLaxb4YFVxR3rGoiVMqvuJkEDZEyFtPVxlGA7sP+S5Zh1QQFeHJNmKLw2WUUh2V9gpj
TST6um4sxUlZYXcfDelZb/D2PZMSxjAYWxog6+XQZbmbBg4inimCZSkAz/CksJE9tNCJPxcsHXB3
GEXMX1+hCKG7sMOOZbVj5M2v0ieOjluNqv4n4yy1cdKYsngXXvTZhZXJlb1ffHL8GgEweIhN7LWQ
fUJEaFcWThTjpIT7+RBD4LPjTocTyWIDuhguH3q4zuckcWyhc75znGwANKjE1VaXStyObqoVHGdA
lyaqtHdgkj/YjZMS1RnBpjXqnbYLNDYUoQh+qflcMCMSFs8rzCVSyBJB20oBImgLpJcW1lqYAIxF
jeofMrvdYWFHjtdfsg6g8SJcpyH6kBE3nR4kzFqLusn3r64jWJW/lM/Klxn7+ePYPHY6LxXdgiyP
Z8FEoeR4NOSgHYTkwVLnQPakt0vOQaE+lyYQUma9LZsottFnc1DxHMyGqBDMHzSxCPPUWJgUo5bI
DCpr6oeE6RMwR3zdzsqsB2V5tLOrVjfH/BJnhomOswWdtvxC7pXUwaNp9+zzMqX47RTqWLjD8RVY
+iaK+LU05hWdADQrNtZAt0FyG7lYNsBUTrWha3jCtJKjTDedN/xRYzD/XRKy2IVlJg+rigV1lnh9
oM1VA20eHCwlPkt6Oqq408sGUGu8cXeHciPUITbE/EAasX/IilqJWRu4g1KXB6/cm/g68NwckWfz
hRrTG8rIOWgrKax/If68jlRGNv7SGZJpimHzfWcRQwZl+/jBvLQvF9Y172VNzkaQZsAQxfClJEqH
h0aK+U9KlrqqitXPygtZKzTDKROBl6xTR5vLLHjJkoj59Gw1pKztb0JMpMSlxdnnjsJzaCHhjHmR
czx1JT02A9rJ8xqxsYMxsVUcKUWL7UVPzmM1eUpyaDGFa/Ixo/ZALofJKc1X+Rj5axB3rHV5MAyj
/akikowWjjsLoWFSuv/fKz415SZf+4l9Oai2dPUi/K3QlnpEpzvA7TW6SHvfn9diayllMq6O8T3t
Ft+J0dCxrLfKi2Ac5V4bioJmR0cIqljdzMIH3DPky6mm+Y3y9CSSdpj+v7q6E3o+r6EjEJWVCSNp
bs8IGcw1Hht8lTdRNScv3fcV8LOFvvkBoB7QpCsrK52Dg/wX+qVFQGNFR4ajgL6SCWYLeAkiza6n
Xo7tqfGy560lsV/9SfCnEj/Cu2K6XoiVqnnTK3cXJzFsM+SYtNmUFxrQc55dy/x6TmVQuhOwYiWh
qtMoUNFkPgfIGJDlQpQYYr3/BRa8j8oWMldzjGPbNxCzpsPu2LHh15TKkC7rFAzgCpoDQ8Q6CnyA
wVhSgJxcSVssAq+H+DRXYONgJrSFlFVOWmtNoQLHJnxgoecaFLz2loDpFW9WG0YW64tUR3hjrhHr
qV59Z7pPJveopfDnMzBFDG3OplS41am3P8L7FX9vqVIQsRW/ygO0sxiMuwe8Nh2XKyit2/HYvecC
4OqWVE3+O99XLCewvRPebyrOW0YoG/BJBMQ3e0Cv3Uwpmma6oowAw6sPd98bR8HvZ2jBZAP/qIyc
hqnXn0kiSzuirP62wI5q2e4BdDm4CidxzJPxuii3eD228DuEA5s+PzDCshZXlBM/O7l2VkXTgq2B
3FcP3J6622+QCfsFepu8dC8EBtKGuSdsJyk8VaeFO4Qozpp/Ij1MBKvO6X0SIfNBSnQFdst4uTOm
MFngru2osCHEFsA10VhPeLL0CKxOUSz+aG2KewZ/1b7v/93SJDOn2gj1kXA6uEa46FQp7LNibBlo
KkqH0v+fq7BWl3o6IWVp/3NNHfXwVc2/qk977Sqdvm9fbuuvb+0LDUJhxEydhHCMrGXCaGaIi66z
psGr1FfHLzfqrqTSDxic5/IagcLJxT9GLQBO1V5oKJv98qkRU8WZejM4PpTDc37Pawa5sSdVVdTo
LEo3CaZi2ynCX0CUkmWz2ehKYmGDQXCsl289o+250ZQdDf8wZX3RmzwgMISZaBL8CUFKtCwvIHVu
JXbqHWhMpKbE/OxrrgSUJt/4wAlSPNlsHBAlCM+FmqrYfLPNV6gW1ivwSac5Hq915p562San8C1/
bEcJgBvNzNFIM8Shkk4qTxzBcvri5EdL/5pBz3eUD80/HOLBZg45X6w0xvRdRSZ5qvto1klg1T0Y
4Z7r/yFxssXy+G6QM1pPe+ZIIMaXTQsTo2joXBqiRJjJBUc5QRm0V/rus6azrUJmmma6so7oCTfk
ONXk502Jhc3JGVJW956YIHsPk4bu0tHzCcMxhYPd+bv0vekEGiy3vIONR6cBNdLkX5y/XOmvEYXn
sudYS7P+gaLoHDZnPA+WQpToo+4cta6bW41w7RUshpY6IKrlD7rKyOYyWIqmIkzpUC1l4hbOxi5G
f1fElgF/7jwQBeoVGgWjqLVWK6Ms+ygeb26nBDyN24vxWqp1eKJfgvD2Sg0xZ/yv+sq8CMLnSriq
Mw9bI2gLyIIOCaBBoO9Cy9g18n2MYBzsNnDWMTj58X/lzRlVvw84Igz8eDmImB/d0JhuX4VIp2/B
iOJaDfUubmvkFC6rPP20kThVjWalLVW+4lu0mvNU8786L3MSxCM2xTP8Yl5xCOs6tUECkjWVfQBv
dAzeSPnTyEWblhcRkhFZI1bbdThjDj50IUmCT3voq6evjOY6mtWeLzwEU5Q2m5Nx7YGU3BYR6Qax
jv/eI7js4T03kmiR6CLwmcx2UTvkzG77toEPpQp0ZxlF7y412KhtAgULsT6EMm8tr/Oqw51N0FdQ
+QQU3xdUAjbHYPtYgRL4ilbBTKf5niXL4WQe53mZQ7Fe1P/fMOy7mGVau01OtZ2bMCYPgzOu08h6
603hTkakI99BSs4rUTJ9H67UUZ0qjuXHaDR32nU3f+uIheyr5ji4tbT2d+S8hOzTHNBojOxKpjGF
WMv8mXobTBg1RaH2HpFeeTwvVb5Ou7hJrDpM0om46UwY4LEhCi67B8tkZBzAMBqp276PvxzEjc3j
bvpu0+b/X4msAfePHvE4hssk3fgi7IgtUe6ctf7z2j3f/hWrXkGkjiEJj0lwoMmUxpsndX1vGaGW
OorruRLJTkSH2hAbhLRYtep3N3rdQSxTmggAhj7f+56rkm6FO7Q3IjT0YgS90yBeQNV3wfg9bjxy
TJNzrmHyzGORBJDpyfZh9xkFD/g0rN/OFu1vvKc8gu/TMLYqVuuozQ1pm2pQXOUup5iTRvhtKICi
Pmdzj/cP31jAzwE+u6r+HA3shrQ13/5llt2Yfb10AwLBlgGNsvrL9ezb/fmX6PDOR1UJ3u6c2Nko
stdYVM3fgLm5TDJc2yMylJ8664+B56mhDeaneFCjCTZdzIuCi2B7WMdffAGMpIF3roFWbhKYpki1
36kPxeEwx1n7aCtDRgOE5DEtKZaUXrKa8wtNPVtZthUJa+6aJYBbYSNLc8+WtyoBZ7zmYGewPALn
5Na9iN1TjS8HH0LzK83JCtWJbZqNv599mEOaQwa2UbyfsCjhUZJ1m19OoWearL+HnPH3g53MV0+d
RGoiSptOMA26LEqFFd9WpHfqsXCB7nZZp0VkwcVoLBC61QpLQnq5YJ3EjRpusHmWnqFOwB00YzVl
OJYBeaHQ5eWIKX8CqTzHP8k4xPXt609FQb5+cFcVgNFnFBIc0jRMZd1s51os4x8yHpcVNOf6bsmj
XtiMuu0T7V9BtftEEwYkpo3Cny89b+odeuuVpFptCbAnEjUxDuSDo13Ic8zYn3ICqtSjRnjkdZ4g
cajoZViVqYxejEAAEEyAjb1AHsd6yXluS0CcN8mLFRTdN7hQeYrVY7DdVvtdCvOjIb03WSQbnHZo
mOiq9CYCvL7i9iRfSehVaZcwSSf33fO/W3LWBvF9vU48CRYJZ7+OamiaQ5FLo9HMTRfU0z6mQNsu
G3H99u29OkJMb1xwP1VrlGS8Iv0/WQ/FBec9ETUilwH5baiBl+pUC2p8hT2iUWi5PvOGSpEvcHE+
Z53ESJE1yHfEiJM5YZMw5EYheai3ctgJ9dsBC0bTMmVrzZXvwF+cf8dmnBJ6vamTB7J1u7cFvjGP
fmsIlvEbNuMDdFOp3ik+hDugLaQI0Ru0rRn8bCWdVNpvoiMAp2kWP7Pz1AGQ4TsHs3N2vLVD/3Pl
15WJS8e4p9daYNhvAEd5VEzIzBO/GkHa5v3QKl7oT/1Olz3O8XcVBKMMo1e3IqYS13Gu68TUIKBa
ySL0OlQqU0dHWfhb8e1GnsPoa6ITWuK52S+Q3ua0oD/tb+/w5MD7CdVfJz8I/MnWghEgziUeiCsr
xNOHNaG2ZHxW3nv7rP2M/e+wn4uTUBYbb1j7kCnblvPfpl2a981rlCoIyXVtO6HBIJjkEu8SI8ba
iO5ZwJYQ51fxeZDCaB8XP88CWkBkzADQpY6+O2KGGr9g3Me26OQpMorigRYd/epixNN5DPsarfei
p+NbGIuh9a7486mtAmTv3C+YuXM+99VlxyjYycLEjBKnE5QABxkniR8NRJyyg84zHVdxEdgs3Qmb
iOjKwkTQczbbEAE0aa71eqqziS+uGyvYa0LN3HSYY97UlUGisjNFa1HfqjEDqrLMq1yQUXFlSGDR
BvhR+8FAlcbqvB+IP+FL//4EJ8D+32tVgKbphLysjyIBdpl6TWDqX1BE9hjPBi13CHEFV38JxPr8
SFXbu2p/1vSKxYYp1D5QYNGrahepkDbXyP/VaRKoL3KyoWob8d5lnNBJlm/2aQuH0UfruTIguwDJ
D10THtLujqk+/9ComwslsaYHA7h8xeXTzbfCFue81rAhAvJ9le4+gKLABjW3yExFMcXV18tVuLkX
U7PAijDYoG3ukbfV1aXhjL+RjOssfC211G4l4pi/xUHF/ags3st2FmuEg0NM6sBJzGJwBgNLCsQv
48zTGqrxWVdhfdFJACZtGA7SgZlLha90IRjwGQttNV613vDFajhyk99uZlyBOiobdwvPHNfc1Lhh
YCSUDiNiYX+r8cf6EiQ3BP306WWU4znJ+EQbWeHwUXajz/vZMqU/rRlcFmE4S2FY280MENbqjsfp
Pcu5/A1sAAhK/yXQp0c5lje/tt/bxqAXwyJWD78MxEY8EzBfgTZ5SvO5mCDj5xY3MEQJRAu6FSLH
m6aeEPr6PswcitaybFXwJfRk3h6AZIBXYV78I/tPYogGPYnBVhBOWgJeRednaMb7AvF6/ZiKyS0J
f38xEczQQ1B96cFnWQPB2LoHcDsEhwSbXnc4IsPT3QwpkV304UPy1sVCP+NvM/oJUQhh3y+plo3M
7RKKOwoLZngaCPdzFuQnmHXX/LGgLtJEJhTWukH8AhEqiS60fJc8w80RGs1X25GQZCUm3CXC8KIv
WWhHGecoLVPk7syFskg0pdbqnemsDAkqgT4lTdlJrYEmYTqx/80riJBBIS8RcU5JTkC7gtevHLEB
fnniGLnWs4+QbJleb5Q2GMPzvNIJjHOv2Q1esmMF4ejTl1VreMNILTEst/5MF7PhXmCST3hLNIQD
1OGgOByGk2KDKlsrAPbGjcQ0uiMLQsiLVWHxObfmzVcPfpdEpvH6zFf/I49M9VD2AVCIKt424LF2
LqYRo6A01Zr9A3a86YCVsGSpD0KCmobHzvH08mIsnJ0E3kwHXgv4mlGpf6OJUGMQW/k00khrXz17
OUnNVWuLyopmErfVCMAdeIr/TGY14iofJ2DxqjavYkYXQb7PkLHC/teK8bmMqW87A5kQHz9SIBjp
V+POwubsg3E0gTe8trdyTw5Qchxrj/sY+EJsxpQYPWITKpAVM8O50m4kXBYkbyTQWUKzd1rwQi9s
FnL3LIzOvtAeJZRteRkpOrDdvgGZlZjQWGIaP0IgIPE7nFsvOYXAcp5DpzfBlOu7Zvt7OOmZ2fYh
K0eOyuck5k+CH0KAXDCsseE2mn7NjHdbNbNK+SKm8gbwC/msL8X9cckIbRppAjxMZ5j7I8j7QR5/
24ighX0ohhHqb7PTqmNPOXVwWssUd0rZb1r3ygUe7AJIPQ+Y3HYuJeRhdrM1VhQsxkXV+6c8d2wo
bfbrGkj7iFO22uK9DxKfamXoXJJcyA3wIewWaSlapE9grqIeeaHjO1he0QJVubDmyJsS0mZiTxXt
xajF3PthO2wWLz2o0hMLIJJwG4Ny0l6MKw2mMlJup3CB9gYaskg+GqYZISXstYJNOOPj4D4pP/r5
j35Omj2vyoHYBWqcV+PfzvbK7pAQjmCPTvN1LEnbQSalbE+ukGtszqOtC17ATgaA7FkPmpS8/mOj
vshawa2jUa54X88+m9XgS+acLohnZy2pXH1gMqhG6qgmOmtq8nWcde9m7/nqTJljMQvDCjg8g3r6
9kVVc9+Ll4voIwYfqGUdqk4AiqUA2J1mx2GiCvznEtsk2QOxePhIiBUPKcZIX6U7YJqjwo0N1KUe
1YbdXgEcYWxspDbTxkMVQpMoKiUXpM0vU+FgGIW1fwoeUB2iGOcSzwcDN0N74XP9eGfSL6F8D9iN
iqCVUJPfeHe0mvFRW2RHOh7vJ7nTptWlfb0jPeZaZz8ZJiuuTTg9fqEO6tf8iH5xJboV+tNq8akJ
Ez/7bIm/kOltIr+sikyC38Ou0EABsA2gnA7PIbHPbcvSWVHHnXMw34DIaIpYXL8k00rQ+n2E6e+2
NeD2eaIsAa+n/+jtz+LWzjQs3ELRzM2BZAl4ZSUHchQR/B8zQuwKvPdf05PjeMQ65CWxppHiaq3G
v6/4vCNeMTCh1DKQWVroiRRNJRdn8SUK0kkPG93/GvckXQk1Ohc9bIFLiluREaGdGN7+ikOnlzkM
1MsPLmeA5hw9WHpBLNOBbycj9x0FRvjQW4MMRX6rxj2B7hdz2X9prbSFM5itgNF3aKhK3m8anchG
syCWeg+WVVYqzNdpxVw0XUwU0Xm30PmnQ8hfK3IhtDNNtfVryF09I3FMVbHgYsD/33UUgFZUpW/T
uWN6JDvCXNbvpCwCwnETAUJW2QPyJH/UmhGB0EpSw6idLmJigiFDV4KzJfR+gh/COrzlHc+rcQrS
7POYxrt8f7bmxDVwTWc56uNoXDqdQHAhmX7xzeWXElXuxBjPhIVxAj47Pjhyk63uNcGhfMIU8OYn
b62ljMVcOHzJEDA+FKq7BdnI4FieyN9mzh0FN8JW2qfp7EOLWx/VddrgWg8NpL0Qst3E+h36xyOT
bRAmush3LhCVXWvyKWfnvcG87HUmRGDua/9rLIec9HbL+Yicj+c6DPb3p8i3Cuupdcag3c84nsiw
1EUOFuUnDY/c4JYeyNVR2VnXeasvqCWPukKIGQ1A93YQAI9LLJxQfa1gGeeT8T+JDaA3mGwlf9Rl
T+Gpvs1XPlL7qOHul+mBRmaZGivsJ14ASf9DbaEzchOqmPZ1G3xIOuNW4+wzCX98+Rf+fr74yumn
xGpbrJWO1Z4gVMvYI0B7enfxY0XrbM0JGusEkeA57xhCuTYEeDzyFzfsjERoKdZlWmL35OROPDVH
iuNXq+tCWGpHn/MYikQCMiUijl9bDD/NtqZlC+UKFXygPY4fHOqgYonKw7Z10FB0d+fRzQ/sNE1l
BmqhMnTLVYB2MofMojXCEW/QdUk76swZIRrhgI672PU2pfYFSn54k/8NeTt7nDBJ+dUInTlBdGBJ
i8iRwNhKQShEHSN6ASpZqggTMwzxmIgnr5I6pnTG1psinpTiU2RsLQKv2Kop9wZx8v2Tlqmy1dzw
iM2ODsoyIocl6ckHLuMRzdm5qNUFqAyHSZRxAWbe5MDtA7rVFXKZHm+QBpTMh1gKkkusisf4Ed4q
z3TnioSpFQtZ0gNkEn8MCNKt6ElJk7PO3LyfGvc7rTDjP2alFy7TZnzNPSlV3CBi9Tuw+Z1tRyDk
A9b9NTWXyVPCMa5o6TEwj28RSRoT83VP+8qioKaZeiQK2HHxcIcAbZMOiPkOeH8+nqIEVuC9+60I
T9DyYXng0lgzqJMrv3eDVFxkxMIhFsfiugGMqSA0PsLZnXOTccwHi1XR46JAjCXvg0wtzH8kdrxb
nTRl5cWPO3dBcenyxQPcLGYtXelzWafxvPGpV+KeVvIQQyvtvFfWNj1S8yi+o8wXm3VqaaRvjhRZ
4MN++O1fxNqfnVLJXBTwE5Fn49nUE/Cjxt9VOD7Wo70HUpG8UVyEVYXU4gVnu4Vc53PN9Rof5b+9
sUDiRk9PgYJMvP8X8mQO+7/T2pnFaAn3S0Qa+5PjENkEIkAOi8hbtYcc1WbkGr0AfA9yGaxtckkv
VLBo/4hk5c4izubV54UjP9FBTxYnqvVVUCxR+Lh8zoepz11lo2utGQb+e8YwajBisGDn9QlrSJtj
q4qcPLcTDygfGcdQ0QOaI7CKEt+VSAKL7aDBqdStmhZIxW+dwjY7j03cT23uhISUyhpn926WshUg
dO0mSe0RWXtvwn6nqFclRtDfXx9Dv+i6kJ0FJK0cREMMicvF2UXHS2vlqQdrHuSJgrm9Id99jnw0
VYKt5gv0XnXmZHLWGF5LhZ/uNtdL7NtylMMf/cHbRihThjW3HdSNSkTAW2f1vub5nFz4ZJ3ansIh
Y0DwyqripnZrKdj7srAAt4ycEyzlckQF0jEcnPzS6jLLdoS3MVfIv0Z05IGA2lZMnV0yE/0sN+zP
+Zx0NP43Eqbgx4rcs2BIfXgHzBwwj/mRb9zBlChVLsHl3ozid2GjOJb1/N7dIGua6O5vincc7BCC
b5HmWDeeymibI+ZUcNAHJr1TykBJaB5Lv6u+SaR01jb9T9rI3lpZfOAGNZmPEld+oVu+xHFff5Tu
OO5diTM+WJwtv+f7WYo0n9YVYUMKsPFHI3ja388ql9nCefTdKI/IC9xwN8Ly5DnOOb3aNILP5t5Q
TAK7Pz2lnrVUKjBO7aZQN701SYujgTlu6oyXNPI1acic1CzyK1zmmhDqRz4Zi68GaFmWfVg1t0Wg
cydVlLnto9BWRyflQlMRYm5Y0zVinUK0k5KkoDFkhxFLn/vtSCvQX0/uFzzdLXXr1DDBDkkbqufk
23NRPYDB24iSSdP1rNM2LKU0sgp1TlQCoucIvWxVNVgS+84RPTmRMoZOohK9xfHdiG5wSYHZb64G
gtUugNbPjwy5LMJ6fnF+IamHRLaeU9luASXcn8EaY7xzUWmtnSyziYVIYpmDno5jlZR8yRmaQtdi
XA3krvRpbIQdZ2nSpdZR0ePKsyemtzxfPDwwEUO3DfPi8Mbwybmn4Vm5Agh8NrMUwTwWZSoKJypk
E18Lz1WNwXBRdieZnVH5BlK4MUMT/5He7TIA+i+6EIUwUWEGGkScJe4yH+Y0jxuE59jAAXUwWp7w
UHQnshWOMNPJ79uKBUl7q4kH7BtnZwOk+R8dqdy/Q/AiVNC9sTCCcX6+xD2GiO9X/Qc88Xjy5EME
1v9NiI5F1Rb614zuOFApCsMTxNVxVjfXUbWbsXyfrUoa2sHLwazwMS7JdIACPfLblQEtfejg5rFP
WTutUrJOyTedmIbQwhmhw6dNHux+zFw38D1cdB09yUhgGGRuP8QGewEtLmXhGKImusYOsW104dlL
ZhNbE7n4pLEmdhgd1q4mAlQxR6VdZksZEKmxZTeR3WCCzijTz0pBUWlWVzmlpvL6MOoSJGo6X4dS
QOcVsxPMqIgMM0XStZuF37Osvre/9sA5gcppvdUuX1Y9iMxNhd+sp7Y/+b3Xtwy/YG1n6JXmxCuW
b+LvRH7kmbxdtceD2wcgos9fyT6BRBvVqW8bWLEGmeNBFXEOasF14BWfxN5HVTERFwnd6bnw5MuL
NSjNPryLKYJMqitYss7BRKAjdIw6qMivIYxT/8VuZukR3WqcfAKS5fuCgp1o7G57n5cwPOhmIknJ
byooj1532pPrbcD/Bh0wSnrVEmkRSnz37iBx/mCTiysTL+TG228WRdqWAiL8OmR/D7KgHqZQTJSw
LXXJ+gSr5qZRhbwrjYiD5t04N6Z82cq3SHk3MJUOnASKHCg1McQNW1OzAxbz5amU5wp99JyZ22nz
lEF5o/zXr7pds8XrVcbL2ds9fQ969Wcc+vF0XWVSdT/8Q/4HeGmMQbwxkqtACJgeV2wyMdn+5D+d
EtJuc7hDGHQ2nAIHzxkzOYoEsSz8JJmr/awx7zzi4YP7Z/TkbieRcKC/LKh2cH4HUnrfzZmOkgPS
3FSQgKduRtmSc6WUrjmsFZBAzPFgf6rEctvoFA9Y9kcqDmiMmygSQHmg7UwNn/SsfFMl8mRKOS16
8BR09fs+qenYLMRSvd0tBf9d183WjZmhQTCNQhHIt4gs4qUev6m+T+tyDwaiIOQllia1Gsc8rBxe
B1eupBl3mMyIEzrjwEKrFTE/J+fkp2Zw2TizYBQhal19oWswSaApXzUsDRPocRvlaqgvTP/G6BiW
pbUda26oU8s0uQ5glecZAnEiNubRrBKgY+7TbQRgq8T/1ed26Pa8f+tUEyjlFP0wnHh2JbDvP0W6
lsw4bx2piqC5t2xPKbTj1X/nwdc3XRuSqf/JRjP7u+2xu0Zjci6m4SAn4l5ja97YZp1p0TDSEsO8
pwabjCSJNK+ktjf/PkJimD6g1l90Uutp/Imd1pK/EeEGboyUDn+HAZYOxE7j6U6DghLVzukWUaXq
hnlJTU0IdQs8xd3peLvrySj1PHotcvc5zx9yIi6/fudtbKwjMs4agcgYitlkrBatVqoynLCyvVPJ
MMK35F6fT8Hk6HeLJJmvqtpz4iTDEzUjfND0G/B3HbeyHa1/iAxg+UF5Ase+XF3eXmP8bD8Hk6Bq
cMg4QKXHp7mgYlgEK1/KepKK0vIGeA9ZBCilf6przp0FqpgMFx32FxXnQVl/hAOAMZle4zXraEeW
mf7zoY3ocfui088/Vp4DBCb+un7ifda4Uzbe6uQmwIB4VRDilBIhEHeUDk2OFGzZWCgDd2yyP6yD
FpVQ5ROMKErmySVfs4FYFL7J7mtBpv0epjSYRFDh72vW2SSm03EGz7dVMw4xkbz4l1WQ2HigPd1i
UIIY9vYeR7g3VySNA8P91OYxmxHxhW7eKiRXtM2+odB1e6Ik2bvIescnYUAl3El2xqqqOLbcmx6F
99rq7FZjYo6KuBzAIrgkvydEecrn/hq1yxnTfNqEOgd6yqurTVCa7VkvWPDibMsSwaANVJC0rI78
XxIt7revI5N4OzZOOT3axVWAVaARd6Sxrwrw+abh6x/WjXiS5srI92sRugXqhII7XyYWrae41IrN
UD1lrAqomd0Gd8wGCipToAuThrfCQnJXqFUToT2pojYw6GhQhZ5OaF1ah7ebraU8/rVpr31GXYuK
hsvOTXK4kUyic3XXIy7Gkae6qOyJwU0TV0oxaEURU/1Fxts6zSyKr/hwyGxHSDn5/HSegIitm4CX
0g2Bc/c2m+ijesjCrXQp/FxEv5cxFeful8hcKHchu1brYZWk9BAaUtKnM2qSQ84ldOsqG7G0Q22S
hWLN6kqrgqqtf7Z22Hvr04QDlQdQI75qFWrme0njVGQLvSD++/HisA2lif3uJLCYxeIhPtgJ0490
+qy52wAB73qmV6lhuuOJ+EnhYMl7EzbWM8VQ49J+3LazF3VZi0hFDomd6fnaB53G10qUajsWi64l
n9HuV4q4KtsJLH4nAZ4WKAOk4kEhmbsYj9vqoIoGow6PC4gTVDY4dN83NX+lW+deYEyqtlsp+ARc
fpx9i2ULgznNHM4vX39uPzU+kfHleWrPeVPUyjcPDNakAlzUtRenzktnaCfW8Pm/tQzN09Mqpubm
YUh/DduoygDUw0crrzi/RYz26+6hMaOGsI5qm3jzLAikBGOCmhIGpv2grbyYvi4MvI68lRZzLXul
LzJIXiLvF4NAXjd+JXDjQvjLOGmbwG7/AR7ezku3K480tVtHTZB81a78EYGerfeROGcLtC+vhjFj
o348WCdyBOgk92lPtD+MfH+TtKhHOXx8zBMeD8YZgL83rz7v1N63QyHC/HD1s/0SCIcVwZHLKct8
+ACSsiBqqf8wVMxkV1efzwraCWTDrhsylvx6hsWLJ0W0E+JF1QKSQLUukl+Y2sGQoHCieAGjXjks
uUmdakLAjS8+6Q0pxlmXHWVRNqNtb+MhsH4YwT3MPKzlQqxKzLebyQ09NhuVhl+Se2NBzWa/cnjR
1A2PHKq51ApDG8pt6918IqQ2SzEBjkLq/mopc2w9/boKx9vRTV04cnWUKORStTcncUequecMxWZc
wXo1ftDHk4bic/4LHcdcaMb5NkOTZBTU9P8Xmis60w/yxYsVUyGQJQBgQsddW/5c3A4DbNDneJUh
wpFASeHGh2rbc38fidVbgv/Q7x3pZIpJ+oA2VvPaU8vtQFRlCohy6qxYbwv3GPxEMryJpawmGkyl
7peOi2wAMv67++q4iO7IVP7hx7Ik3sqL8nEs2Q/zyO2QFULEQTcepRLzjRc0s4gbDoUU9K6NQVQF
bO4TAgkJjfRixcB0zfZ0UkKTX5QiuDs0PillgiIMfssYSWSTAOjfi0np4pY2ogge60MhOMwOjq2Q
ON1Bz6rqmfEOK4/ptmuQYxBMFuQWIDToDfsBV/y+mPQSqk8eM/WldWfCiQnf27pKZuGU/LxxZrG8
n9IL+vUhebMtl6ce7t5s1/51NXJmbyjpjjlMpXNlFA505yGdpTPjH2hiiDIdQc0LNq1LZITLrzMZ
Roj+hoVlFG5ZgbuKaBK4BhoDmGiyLGmsdVVu6vU9gqWVZPTatwud2UlDP01tVg6ZKlJy8H9GTnbt
eh+fcVGz4+rGzmcVf6UgziBgIceBvESlwC7xVOOFPXjPU2SH0sMRvlnd6NsO3FMHKW7epcwv0WVD
vtFbQgvUhurlewW0Wxq1gb7VpW615V77oweAvgltX85mE7DxA2Ivj2QYjFOPmRK8MYkWQR2rjru1
f/ULZK86P0p7kW/YkPp1+sav6+nzezcnCUrTjdAbU49gJXn8rkbkWeOngLJA9mUAQLa9vrt2iWxj
7Za5nNln/Pe/ggHDzWF0bj8UhFZBP1ZYAMg92RpTjGJA426UmB58UnC11nOtvbkLHhh4h+UFgzDH
zD9SbYCug6UO9mku1/EY6fmdTdBT7e7nRJtXtCQp2AHNiBwCF/pb/v/sCnIuA/a9oX0vay2UE1rl
z+C4A0cwQbujUi0Qm3uNjjq5zzBQT8L9UR35+Kl72XMLTQ+dIhy6owuwdCMeeqrLM9N8txIIYIEI
LURB2s10PJ6Gv7tm1QcKSXvc2mFIEKkfIBvWrswDF7EzOKdfgBc90yydHr/YJNW2RzzDd+hiGs1P
vPoj8P+t/E4rFd5JZRAWRpjhcy9NYsmN9ZBGFinmBpKUgcc42jdUyO7DfS6eBDPop6rHZPj5fUmT
CIItSQJkulw/gi3ELWCKcUGlXfSopjzk3UJagAyZFNgymAl+4hAQ05LV9j7N1zHAmfivI7J4y9lh
D13YmeS+L4aM0XsG+zdVaoNX3iSX+cSvNubcSapTjnsUOauhqhr7wB7VD4R3pVOkNmrwFHW2mFcp
rsJI56vFYZg0L/jVV2Hdd4VCznpzGEYLaIVMegyPQ94essH0xAFLxCwVyzYsdyme2reeGlncNAvu
OP+2fA/2rgYWSAiij3OsSqVBCyEJPXN5OTDqJdAUatnUcJIcwzSeRBX3RN8qcAJhqIosDxuGXwxY
qvqOYNvlGt2OGG3bU9iYojAd3mz8lOksVE/OWGt6u/wXDQEzGx87sCHcWp0yYYqoBuv+l3rmwveW
Dg5t37QZlgq9n77cduPiQBtB976/jfTumSmpAGxnoayGd0cQ9qP4Yprs4C8uoZ4H4bfGcqJdZaz2
IgJMk/GUHwrEJcCtDx1MV4YpMCW2eO8PK+w0PuX49TP+a9WRVyrERyhW+/o0PdUryoaN+XUpxl2k
fj0sG7rF+Hi6RvNbR6RiX3GiWTGquMRZjyXg61/DwlV0FAcz07fIh/s5HSMGx9IosHiT9PpYA5P1
J9N6oKAqt1uc3toxLVmymx2dIWYvi8Vp66xaApya6S/CHYYCuhSGdm2HnasnQPOioGo3fAih43Hs
zq5j04l15geADTyruWaKJ32Mh+bXFwj85Yab3KFN7ln85Ahdbc8jskaA7CkUi1UjtyglNv9K8iCA
2Knw9AR2gsD0++/wbL++ci1TCVSAHOzUzWdlYN9VYDGjX0mHWNj6sE00327wRazrNQnPmiAVmys+
RTLzI66TEmsuh02KrRDRwCnz3hnQihUgjBLb5wjuRcV1JvqpR4+gyDBtZpnO/JwSPPUD7bfqyrOo
dyXN8VZYX91ZR1P53YYIY6EgWo1ZVYnK9CAYFYjX5ah2bOz1z++yVDj092asuk51FtyemtpfFCUQ
l9z0JzS/aBULvgFNYV/bCtl+h+3iz8LFve/vS8VZbTSQLuhmoXDfwWu+U8Q3JzHgXArDjRMJwk8r
9u4RmohPVCLw9DZaC0/sCWJbzqItr5kEnLRa5Y580sLOVMoi/iOOUzILHN9fDtqIHgmEvQ/pp90E
F3hKIH/DiFQIDlvSR4+IGFaP5UUoGM9fAlxqTQQvNHSSR78pBncfr6Kmy+vOe8haBWhDWsDXtDn8
yehqIfXe85YBS9pteZ8hrzapfAGY59pBlYLfejPsqOQn/F6Pzi/MoGZPxEZFeNGiuh6GLeVXn3iF
Z2Fj2SFcCJHZTFLdkUnUNEk+GBAqoKO5SfubdYbQaX40mWGWmy4xp98Gt2i2ZWswhqYojQU+mH2D
e1j8Dl1big7f6Psnopw98kUCNYL3KbU5UitXHdHt82JKuhAD1GaOKKO0Qn0bTBNb8FDwLSjWjyHi
ssx8dyDPJx+AN5h3uKpnKfqeFlVhKy3t2h2krKoSe5hUqlTNtA5V2BKH/331QaApFn9EFvh3dz31
Wc+VDzcpwhYpFaVhAks4Sg5Rv4UaB10M6PySZ7T7SJlLLgDyy8u1gaxkh3fc9JBivLIaueEPOB7t
m9oYYmEfA13cQcQkqxiC/HWIpcJO3ACfWsvm1rFlwmT1gr/df/8McIRlpRdUW7PPfY35IDV+dan4
uOvzhjiksz+I3H7nfUfA4le1WY6w3ijPVy4f7n0TRwLrmgzUJhiXC4gBs+2Gk6vZabcqMFH5dTDY
as9AcfmFjUblGTAfFPCmLX5wty04woqyVo5ScPkmM5F3XkT7YQSXS9P2hQIhGnpRzy8g4Fbttdww
2oJMikqNpKcnHN0WtgGkA6mLnLi6xK40Q9bxm35utbxdZlkZM1wAVtmByjg/4Rpnmdbl0pLXSEB9
i0X+/8rGqlIGvndEY5Sre0iihwa7Ae0Qm/z0R98NDPXWV/FwptbLUSYOWATn5Nu9auXb6CK2tKIa
reHXAqVlmxLdE18m+yH9iJnpamhP/TtDQpfTKqg3OCgPp3LFGea+t1KsPHSeynWT19/39ytUZ9JU
rNhRUtbP3bzOvw96gUGJut+dUP5tdxrzwhO6duY9c+uyLiEICvQffUze+KXY2XBkEOi8uUmwbsA9
Q7iLP1LH/LuFM+hDJIwBg+62wxdhcq48KeBvJPTePRV7TFR8WHguEVSo9bDRXA//cSl4V/L1TAS8
AnY2skaB0orynytJWwWvchwWVusxBPDrHg9AbZI+DqEAENx6oguzttVky2qL/ICqR/KJooUkT7S7
wS9LV78j8socn+zRmgEwcWo+72dSJgm5WDtvIpSuLYF0eVbVmVzZ8mV92xnAGYhDHJyfIJWuQutO
TaAn+IH1EPHRX6VywXOTVo2e7xkgJekE+MMp3PMy9hRhBCkoJi07d+O6rE7rwsHqCVzVkDfbZLaS
PSiZBhL61JdBMY90h9KggguKmfBcm9TKeQQvFgiF559G0exfp6d/DVTUolmWit009j+YZF6pG9qw
1K3BUUUYs1h4brx3dsNx6/jSyEiAER8d/xNKFYxnqmqncOmvKfLi0U11E7ZMVFBm7VudWpC01yta
WNIy3ky/qGn46oF9mPxzPzAMYfqXm4jJeCR3zLgHx6VUV4ZNLClmstjQIwL3bty1BBmvZJxXYJ6V
zzGYACQ2FIdgvjJtynQyNonSqDzzACQuPadQp8qtYoO4rPOaQtJJa0FRMBr0R+u3Q3x3OVyHHXiX
G0GzUPRVjp1hsvJwG50D6dDCZl2XL6nZU1Rw0Ob//sBvpU+nYestjG/pugZEM8XlzcZcq5fF0fWh
u0Lf9f4pE7Yf7ZYQN53jM7SNbSXQs5ZvjjtARLyuD5gPJXjWge+32ICo6exNZ6ZXdk2uvB3KWy3X
jSumjTXCk7wUd8TZCZmynlP/0pFf+xhVYzGCgf2HxgdPl+7Bl2S/urBQlgOYs+scguo+gJe4YZ+B
1rEMuME2lLXBLvuBHInm2fpn8ezARqJDkxu1vV9wGDg7i+NW5cYIPw9bnzgWL2S2Szhx4V+qmF8e
iX6fQA1y+LXFPtae7m09iJTE9VloRi270ULXaS1oO8A+OyYCVJRq2hVTRBClIisS1/8E9zLs4fph
4mCrZn8PXFwawdz3+YMZ6txPG3cMGTIwoWKpwsdxaseHuQWdUwtzLPUcovyoVDyZB6gmtoINXnuV
KMsA4mltz0eoGiYdXMscezGOw8JrkZfU+1164n4eyrLm/61mS3udfHQqJG4ZXSki0eiFwu3mcn3e
1Tmootw1XGapAoOtUq/sKv08Y+uIYg1J60fk6WSLLEAY6DfFHpDnFBRYx5q0f1qjIhwBVub7ZW9K
vbtyMV1RGzIwVtxk7Rd2XjhNECkHaB3mwsIQdNMJnY+BgMxqKfNilDVdq77mbCT8pN0iekpiF5Wm
j8uhM0ZrMlYVCEt4RVVzfxM1KkEY8N6sEcy8M5uKjRdQVjGeQagpc3/SSV1l5sXtMp9MuJUwHIur
Hr8Lun0O4v0qK6tDNRxkKEo5Inm3jhg4+DLEMeXFB6IhkA4xmQF6/Yj4owciihOuHAA533GC0b0E
S/I5Pkn+PisJDu3OWhn7NZ59l0or0KdlE3CJQSijFhVazvWxwOis9DgOkfmieDx5gaH8d7oHdz/R
OeaP0vGS/STYN0QkwHClTBKEuIRMUViMKEQIAR5x9IIO8gatz/4lr0XDppuTvPTURPtuecSn2pq1
iKpyRkRfupD6hvulo9D3okaqFToW2awDdg+3LHQi3urp5jxBQzvjLvWocf9oCVjp1Z+riSi+kvVv
l852SGlEBS4B3MCLQamrduIYuo/OsXLh4Lxf+ZbTR9U5fZMgUvdEtRBdFEtRtU4sUaHaJDr+Co1N
vNiQc0Z26elJeEPtFa8iOxxDiV+5EZhe5zjiZE7q23K/GwjynOoVYO24HYZ+NdwHY/jpgTb5AaYh
f6QRqsVzWWELIey4xSZ/htqTU8QzKC/N+y3ofruxUN0AiRojXwr+gM06ePU7NWJ/TerldSPanxCr
PsLRhqiSnqcnkRK+xxPXFQ0OMXU4Kpw3dHHqBDF/HbSFtzh0maA9hJnIej7ri78Mhm93IvI2MkZU
WuDL4pfbIig58mEVVP1UV6gpJ95jvdNbeOfRbp41V0hSe7tRP573PjOlCL+KsdOVAW9rh++BLWz8
ET62O+RMW2yPEOfJgcKfDj1L3dM2YpfAt2fTRV1q/QTWbYW+EfejCNBUK4IoHom4WRoixZWis/lE
uNGKFcAUSXvYPAlBFGBEShxmsxesVI6Q6ljGLiNwn7WqE80F0mjXDmQ+YMRdwZx8sj963Flw/FHl
WTB3+B1DPKE7kE3GfYWogFvWvS6tgIaKWGy0etnbSSK9YIP/QZPgP99Ms0JIEPCuJDW+q2uzpZBM
C2HsCjbkRrxt2dl+cwzG2BdQMpIHoK9ihWFZsQqlx9kpj2u363NKrVzbU7PvX02rVWtpq+MBjD3A
zizbNMNlZO7tAd08DyJZM5ZiLvWPm6EoE7eBaadgTSQpLa51ZwPt1h6+t4zQVFIo9scPpuQJ04Bt
ya8FJVtOAV6W16XtVnXjhKnrS4HXcpiu2DstRyEFthAnlp5RZ8duU/F2+R84gspjeYRyQ0kvJRoW
wCimDW/NtmG4Rh3xBDWRUncU36DWLr9Z36elqTiIqt3gCgpKvZwWg+lRLvHwEmc9kiDfsXhzWWhs
IiFYPhqqz8Wv0LG31MOrxEdqO3LNMrPPRF1Ug7WfKpYQj/x6bnsGDPMkw9WUIpRnq9NT41Xt5J7a
EFolcgQDHZi7RC93lfzkovVHLGFT4hDdq46PEVWfMffwr+TuVQ0QEtTRL3Z6Dbm2/ysNHnGyW89/
gbzKOMPNKXAHt9OFqUuFKFUoJldU5IwhgBHWqctP18yUBlHB1ZVAlLvKTPTmsCQmkaratSXbTOQ1
y+uQCVm7VTqgSKqgphxGqifkDnAW5ax22S511KcNdeSSBjTH/dbXqMw1YucYbxTsPd0yXb/VCAe0
A/s8r5IJsklsa9sad5ayziSoSUZQkX+6/Noaqzi3ffZOPuvvyyOrXxDmdHxvfZ5zikn8Vu5csdnD
jmFujetG9Cvy0/WNaWxgXSuPlkZjIIsOK+R/tBpV1VsKbWyQjY7lFNHIb8A96/tXMoYo97TL21A+
oB+zRIVZr2M0tGaCo7D39wdaXdQmFOZfMLDupaJiRgc+/kRpLBN2D0U3LJMUDJlKQY/fe/yimZ9y
sfExLqv68dEn21LlsMQlpgOjb/KSt/byn4LegA6u8mwS+ZQojKVmzHhSb64Ka4p7VG+bLR23HfAH
MGytuJoS4M9zCMvSPJEWEwpx+HiNHzmvzrPnXAFw6idGDhtzOmoaMjFptFGUuChN1Dqxor+TKKqt
de0OFOHBLXpOM18Cxmfeeje0nG9xjMARCncccbVQ+lCPbhpcd2DGA7YYwfj1ubezfS34YVP4GZbt
59DC/YZdm4Xy7QAIi29Ol9J0P67+Omy+Zb2c/9hZhrJxgbt89wRCpx/YygYsdz1lCSvFItqeQoet
d6MQ2pEDAcZnpcUJY7wqsHRNdU5cgNZimgiX7rMC4A2kM5VzRRI41CPodb9iixQZKwnVGsRW7yAy
N/R3gRqISRu0tRYDS1+ougTU/0M98OCirjwacMg2Z7as0jtuSEnLxarcVERwGf9f2HSRIYYMGp23
SLm1szbRRGJ075EM6i2U6G4gs520J855lyhMm8Rf67pSJaQxpRFd3yFpzOtqwi0uMwknGfICIJAE
QBZWiEThuSrCjOr9duTWgTg6gsRIpVkR+vfOaxTbL/T084j1kNYjoDRHdXdQa0+WNqbKawUpacez
WSbEzJH9q1IX6dQ9Rp+V6236RKkJt84C6u0BBpC8tjHQfytZ7zxD7vtvBEt6fbQtkofYrVUfNUom
5kfxloE8H2H9KpO/vYmLALWCnuhTLYya4nSojbSHJsCUF/d8mYT726oGTEFmXA7fRGElJ7Umshgb
VyvaafZJohkQxrAUBfvJJv434lRCH5NiseqNej5R1NmJZ8NaYZOAlzZlC3pXXvDmRYvKvNB2P15A
yxKD9i8V1Yoy42/4Fy66Kghsfgmx4q5SDcg4xqqIDfVlMZ1jLdC83G1vV4ltvtptIhQszvQeOik0
rTccCBw/ivnpp+7IHXYHbZ5XhbIHujptz4Dz8RMUHr7lujKWOVKyQn0kSMF9ZPXHXquIQd+lTAyE
n8jPbb0GxQ4Vv7/O4TmpseBzgYyiddigWR/HTex61tLxYHiNCIQNetv5r+hgk5r1niZRZSaqDlfC
owGo+tqlYcmzPPat3Pvf/9ZG3FkisAFYqm4h53c5XUD5zgd7qvaCROQQpq/xRMLyAfr2jzhHE+tk
ZuSjF3N/sdHIFc7KkNIW1cb156ohcsChxdfArlFOkRQFAq6pwo0I9zQdwjM9ZcFbUyHZzn5gql3w
sC81PJWMvn7aSG2sj7IDwKBZqhaTls/ZYRHgiof5Fo0goviqko0FeGadlTySxotRzBCNjTUIv1em
jRaD+7OPFmuy0cJxghHfxfUDJdQ5Lq+GlQy48Sfaq+h5zed/8w1he8n4CM3phkAldoQrifoniPYa
UIyk0/6BLcyDRTTXgGqerKvzh3pCdjwqIvVanEuno3oBM68bWpZ8ZkV8/gqUuNbSJQT0y7qODR/P
6XFUeHjPzsax8ItN+u7a/MMfq9WO0JF3+glnBO754xM6Uh71QwL7d9kdiPUZGLXJUjGo8SEhv+q7
slBNIGOGHVZjo+C+hvasR22BbOKc3o7U90tGO4eUz/4RnmdWQTutQSwNJpjzS08LY2SmANIqA861
lgE9jhBR0bgCib0qRbJEW4KgztApbbItW3eF8GjXp1HwnPiloUpFmJjCY6J0BJXgak/gK8VHpvUh
w3USmJc1v4oOVLuq1qBnVtLNJtwGgH/4roK1dBgFjRllGLbR4tcdlbKpr/8lVRG1riCIc9VPvwqi
NhXT+8lmk1yKvIhTHavkcKcr07r0oqDZeozjtc2cREf23CC9DWyX9Zz6x1+2fvI4zgE8ZK/tWZLF
DloEDYJwEYja2Ncg8hbQCYh+1xLeplYKmvQDMSO9R5V6V1SycsIjYU1shTGjesSkCPUrYHKh/5I5
O8tJ8s2mvz64KPwk47gYsqpMCoIgl/UeZ2K9US6f1CVG0Y+PaL1Bz6Rl9omKM7eJDEVEj9SP73Tg
s96hjdH+mkJC1ZYYJHBAVsMJsbbfdURnB/S8myc8qCKCHjDCUi4mg6QoFGIDLa6rxMQRsuIqgI9P
vas9H9fbwBMIuqE74BJyHxeU+LU9XEt7YfWTcmPJv+E9fbcWGIqe9OGVHCwgKYWdOPOpNNCdG2Fz
KCVXi6pjudDTMfUkQBRqMMbdSTkfxxhVokUA9B6AyHVp1ewsMYVSxjfiSQWJC++qruo9ZTJ+7z5P
iQbuyoxa+HBOR2xtRKk+MBzONBZRSVOl0dSqX6vBap7hkzbn169IAcMDlX9RG5MpMllen5KHN0Jb
WPv2CKncsk9VU8n2ELJrBwQWlqy5G/HELskXtBEFyGYg3vQ1AbARTv9Hrm4f3buhEIQdzrDJBkU8
swGXeFqcFfGOhQ9awvxlS5e4GpEy6fFnSF8mk1DmpNzeIxJpAFLWgvkoym2U64TgHlYOOdDc/w/4
g2T31tp68fr+CLAETp708jbM1+i75xWPPEwac4codDi8z7WzwoitZhRWytIi2lR6hpktb8JQ/iwy
NVZY6cQoJR99CyYiwCyYwznKwUoF9SMjY1gvOfbTLKKqQMxU8s2A/Tpp0J/yitvVJt8jceLaKdWA
Nakv2l704hi0O8cMHiQATiONR6BaSx4nHMlOkWaLyk85jzk9HSVj246tPKCZGyymV3LEr6idXnqt
rOAYeGH6fXWPeRfuHGKdtT+ww2gbMZCJuAzPbTdxAFV1N0lS9sTktLnHuKBm44bxm+g3i2165bnk
u2gcVd387S+za9j9EFDe2A81cMAcmANFmg+ly4dxhnH7MrLJ9GPH6Bj1ld1rAGHuhnZv0lanzdjG
6G3x/POdSjMJwqsRqXtyMSC3FT4XDwAGXh7KjXpy6b+QLSzaN/rRYWe0wYYFL/mDkkRiqiGYsRWx
XYJVyDq9e+gYSQ4Ib84XOBX3FgG4TpV9HtXZ/18XugZILHg4omozaEgFVRm/5OLj7paT7AekUuxG
AYnxFROdaFYGEL5raMWmV5If/zqO751mjKpaNb1AkZW6d8i3BreUSfGcX4+FuMeVo6z4q0vOX9xt
QLpLkOtsHnagyuSSoyfY8tSZBuChrHins1SPGs+HZ5zgJ1zfnwMSGlcvWZsmB7qOW3tqD7yFBiTN
f5eQMMC/at090Ye3Ja7KNbboF7++vvau2O/EsvlaVbLWUS4wbwIJvJsPo/QUv2pijPahUafppE+V
daxpHdGEyraFAKPTVC700uB5EWkvnhx1vznBVXWblxGU2DvQ5a0hjvPBs4wG0h8mf2htlM3lo2to
y51ASD/6V7YEX28hil/scg3blWvbfd6A1+xuHVTAE3UbvKkyKDQRYXfQkUhy60xpLkA6lFZL9Cia
7B1DmF1DAF6owGhf4cOmCt/9cdTiS4Rlvuwz7cN6wlutLBoRtuQvBbJkljT6Ob6bSvDCpE38N4Cd
cxR9Psw4BCyH1u+aeoyBz0SqsNJJRGautJaj06UYzuhz18wudeA6kwdYa6K7FmNnVb0Q/ePYpYNY
+dqtvx9OK/Uqj4N2b2fZQaLtGt8wGWRZLumKYk+HdgOI8KyE1opdTghuwk6b65b+597371IhlSSR
9sB4YcXNHd+/50o34mF1RI4/NySeKvm6MppyLNOSE98me1r8YmQ7i4RMwXzDGfC1EhXH/9t2p5+Q
wLRQTbSn3pwunjvDBodPdi0lRfxbjLvDv7W7h9h5AvpZO4nqyj+UXXuO7qCEBylBJwyRmBdK4Mxb
HqqA7FXs9nlT9SC/gdqj04bRUIVDZIV+rgGGsMEYjExPYksETNwdM4sgdu1jV3DyyP/6PqZigTzn
8b5sJLJhsgmA/uDjtQnAqkbp6kSiaWsHc9B1DoBn4pN/KJX65tZYOvx+jKs43s49H+D4bTYwgrnw
dUq5Tle/QB9Oim+UJbMA0ZSrsgkFK7TSutaval0cdCeITtPTGBIoczZTyHNVHeFF5NjXXPJuCGN0
0ryWo8W6UeZTeCVwKXnjOfq+K9VyPDgGf1ncJsrMmtMuIRahMrVtwRVZXOEWqyFvCwy60r9VN20j
1FfNsc3Uh0YyMqBDtwYTl3d2lMICNg+DPfMWNDroZPhtFcT4iXiWXEqFa7FhSQlgRNW21sJHhhuq
fMpzs7KFVVfVuE2q01bU+Dzdh3ox+TussbBo0yzU63UOaI8swwsdFM9JfzAH+GujmitOqOl51LYp
7xv86HhpUXlr0wy20zRR8aWmQbSyeP/vnnq0RSBhUWoMeZOhUiy/HNNlT4K0H8dDuxChWGreNHy9
oXfTSoxYQy1sYaC1ZaFnbuGn/dpgxlbIqlQjLuzRF0+Iw4NnrbZmFN9U7FhBVuO4BCFoZYu0nxVI
KCCfSk2PfF1LSukhEPV/qZ+BGgCybGqxUJlLIRiRU6bVCJz5Lhtq+eMurC5WxvEGOA0eyCnXnEXy
1Ti9B/I2GEmqcy85pMjqCjUlU1/7PqWCE/xxiRN1fZAPPJiuMEpVLmQyTELoGdB/GBeLL/IQEtrk
MLqcjk/FoyKUkjQtjqk5gKRieZO6LCNG3LehRxof/O2eBE2Y+pyUNgzIvetVEEREJzgCQgi+7tN6
AmBM+xaqWasiUmyLIFkgzZdt8MFHq/3U4q2LL7csKP5eUfEmHOkMSscFg2ZvqY2BAlUcUWdzeoqI
ljWTv1jc68fH8ZVPXiojhZZIcX3ztWXhklqzIszoXB39jj/Bb6kZ+feYWNeb6WOGPAQKY89b5ZfX
QV1h1k+r/QnpEw+6yNfKiE/+bKc1QGtZD4wwwNRlsWeN4IstyPPeQXdFwEJZ8gv1Vr4c1G3bbgs4
jVNIfCDKR2+eBZme/DxP2Mtot7ln+8NBw3z/AVAf/HBgNaxgoF4pnNXZV77s3GIf3sqZLKa4zt3i
H0q2wARDTTsgoYN804Xw+8keAg2Z4sju5twvjwR2xVQHMXB05U0b2CtV0I7NDUao43JDzw4ZvmKR
1XMPLBCEYDhk5oncgKPFvIE/gdw/l1+wonVaOlGGnnxJZr1UoytzLR4rVTUTtXu0qcd1jApwN0Lx
qvT1kg2Zq1miqyA1Cn1jts7F5xR6DKLzyDZcxwO0esv/MfRSkXxLjtp+AWTS981R1YJEKbvy5/NU
p7VjfBDqxohtCb2x7/YqKX41uPmdvH2mztYwds4pJA529Rw2z2H+R1NEnLVCOoSE251mdk+C1j1Q
0b4wIzNZ7cBTA6d43bni4rWhBpyPI7XzHSf7wRur49qet+kyuzJVcl5BICAKKGyyvsjQTFRuxk+P
xA+Lzx1jkIznO90mV11zJa1lv1qfNkaia7b2naWf+FbpVuL48b2EfWEYchRyFW9oPR/VcNE1K3Xt
tvznZVjeWUZfHjDTncL5mDuyRDVRCP0+5pj0Qpz6auyfUfh2d1WuOVkYlf6zIOpToyP55Y8ZxRfB
RS70WTQgfBAuB2UZ5a4DAYR10qsbSJXVKk+V00FgQeCJehCIex8LAgo0/cKCqdKetu0/IEa7HKLt
2FTbiHch/QhRAA2YcDa0i+/ChlaOe898nQkfOENOiwLoSG96CrokA7CXcHiGSPuh3sNBcdrbfUuH
IDutXO0ikXT2rGE6Q2gafy5gqr1eVvtTkzoRBluSiLZW4HQfBA+ZHGm4apfDrq1Io1fvzEoLCEEa
/w1+CaZq2aJCw7fBBZvHP6gqQgoKZjQjfVlwTPGz6kor1f7vB6zi+urX9dEpjrtpP7Y+kPChWv9i
HjXx20X6MOs39YQzPQVScP6mBqYXKb/T67T66CnYXEsz0YySbwTYtgjsEJ1gOsSu9RtMZTjO4OuC
yQftdtTGB6sgJF6qPwHJRNffX71pDazAbFgTodOC41cezZ4oJrLBWlGaTQsYaFc6cH9ZzQccbIyt
7xBcTlCeZdqa0SkSgs62YuRZ5ATz91t5x5fcWQa9YAl0w+X0F2VFdT2vggsbRDr7fmNBI1FYkpHr
hS4LoDj8w7iAVqEs2Y5TO08cUY9WbX5EnH5sDYMvaZLYDxY0kTOWK01WhwOSpxcg4JkkBhPJpCSE
F1xakCdOU/ISsfcgCFZ1Q1lFy6Yq3w1GOmqtT9CNR1qFs4+qqHjFEDHule0/an1R54B7NTqTOE/D
hIrMEGzBrkMVsZWd2Eu6n0CJD3YDEyzkRb0xgOSswPLTR+TosYvPKRGh0TqZFuc0brFyC0Cw26mU
ZglXWumiV9ykUSiqu6A5x/Ja+5YAva95nwcqiTeCQX9hG7Dwq7/1z+5w8G0OsNhf4LjH9fXpFdA1
CN43FNHlbFACCpXWQFwYA+eJCMZUMZLmTJms0K7rT2fgjm9SlKmARzqgwAyum5yuLC7rz7G98Gw6
PQlHyKgXmoATI16y4VUkGaamKVlPO71qaqgBHVp0d+D31zrOVRplvczX6bl5XLjH23kfMOS9E2Qw
iqAkiD4cyceGAtq+TLufybMAz4prBz+Iq0fJRhyDq+tZUXj/1uhzppmbC1uqgKEpQBnFmiFCHNDh
W77Gz3ehOH/g35WTavsQnOa8ESnGJWCb/8GOo1EmoyZ9fbZuxfSur+QxsusMj4GWN6HRax9+xTCi
Y046+Bq+H44KKiLf66Af9HmotiPVQVSNHmiXqdklrHmzqgEMO2xtqvo63ApgaqRDKa8pHT9N1kXQ
2Vc5JVn/spZE6ijQ8e+Y14e8B2iPkmG/WtQA7yDq7qe2UVCnRGlw0by/H82Aa/v004ya3QqvUluy
4NF+sj4x15EYBeaJL4wy1WniGw8rlkSqs6kvC7rTlQDVfUmMNOano6ZYi/tpLbK6LsBn9UZgwx96
dtW33kkYY7zYOBxDU1mVTO/NOKVGtVMF9ekCjc1pI7yckf5UhdT3B+E68vhwL3KtT3dO4cQh9S53
zBbZOAvga+hF+PnGnRx9lEt111AOT7JX4sscliWcSVQ5Y+s9NOXKxJK3JZvXEzOACDi3px0wVVOT
WUWoFjcsMGG5FX7iBQldtTi8L1qWd1v53B9/4Q7eHkO+9A/gtaXgHljFeRDw3e13P2mRo5bfqqBi
qXWCLMeMFRj/ZTwUjHJ2b7bI9kpo8ubZ+477Sa9NOZuZS01IP4/azsls35MeUVKgaQ7SCPGorZfq
C6k5M4kbsOR4gS+10Pp4DW4Mgt927J616HPqCOAGhb9yffZAWfcd9L1WVDq8qE0abvogDzENU3XN
Jl0WRm9N347Jb8nr2D9xdfceNnK9dX1HiNGniPe0WGswR4d0blU+00zxjmVRleWnyQ4Lg2guXeTS
URE3VpSkg3maGxRtcxKBcRYgqs2YQDHCyam1agmO5V8kD1br7a7NlEj5LTTk3NyeuIRvnFWFQK2B
ZZI/dMrsdLUyJdZBCPVQE24a1EzNHUxLrPd7w7TZL4SfShT7KHtsENeu3efgdMUGAjvDJwsfDHcL
LAU9JnLYF6yeSQe71d91d24dcKopGcylA1yEaNHnAJEdWA+LkQiYcfMEeAa1zRIK4W9LplrNRVnY
LVp+HFdvLZ3F9FZbDUFqYnBUcAOOR02tsWYIP2/aPZBf2aWK8DV9SycTQMZx2onYLHKDa8JbWmzQ
ga0EeJqaKYLxng3a7cNE/7StAx76hfmgXtZN5lbyPT1RKcwkFzBUyptaFapJV86twh1aonlE58up
MlNkZoSvlmnnXQ9AoO7n3Hue+TcMUMTTU6aJWMkGmZznQEpBrQPeJL7eclv5spZYxYs+D9Ee3tTW
dnD/Olh8++eVzOgSfWcrtEyoX+V1zkNB4Ce9bwbPgSLqFqnZkOnKIr04EPa0O+lvEy+CISx0TDX7
QcKz8O2DkNEqRwonoPYJI+ekb6BvAK8U9ziCtTuIYN59ofPUFYk9WcVbLRkXqPlj7P7hYX2WJbQv
2zHYG5ez+ui6jUzTOzMb6ExOW9XmyGESBFzPUTjHbWhCAJaHNJpstXCXhCR2gnk/OImzP3UjM/Uk
G5uKuqnPSN3NTB8rlAKEUXYOmw/SHIa5HMApoMoBDwb2vbQ8uXX3ap8s6DaIzIhfwnZREDSsrbpk
GMSfJXavjQwg6anMAndJaFkM9TT0RkSBDSjZOGo77++y+5g/fSE6U5ZEEYvzFqjS63RV+tIT//69
3xYG1dEwk5dW9wFU6ChIBWbx0iqjMurXL++D6f4Ym6b6yRL5RiYwttZ5TQICoHJhJKBsLyeY/K4n
f7L55VUGtwWAD9FJXLPUZhRPu8Tu7A7yHBVcdXrvwi/hHHCps9F7CZ7ZiYxODeF+1PWFnSxGV1Rs
Q6ZQ9R07rCwpiPYdSVGIF3gXm7sKdzQNNtt+3TvIHCxuMpLnMZ7qN7ISKGDKDf7pdpl60j+llOLf
sK0THoGxxyE/Aa63YGNNiNUJsZJD48gk+nYZc6bBwF5K+/sF798F/zUWIU3vngQ1iSCzZHmlbfB6
GKCz/6rczpptSWEeIOY2v/6TrSk5jY2vn4PBrJrQrdjklXlLPM/Wbpmdp6shwSTJIjVk+G4fCBlQ
pzB5bbPIkbOF0RBm3eeqEyvH6Me0RS3OQt/Pq++Q0HyYvRL3wO+ll1wQfHiWn1ZPFHwrFHm7nHNm
yx2w91P0iedGoROt1WMc0/Aa8Ag7Wpaq5poe7L1iQbUqCaxADJxXF7oyIeInPIsLC+FGr0Jn2+Ix
/i126q277LQzMKMksvv11lqdTnXXA+X1H0UmeLgh1Qw+AThYBl/qelc7GId/GxPdwDRYijxhMYxg
J6CWURvQ75bclafqktzYHAYhouei/uFhZ+OFnwS6MmFae6eKy3RPC2j98Cahct9hOfjwtkj+Bsh8
GVgu4F9LcoD5zAmyoONFBMg2TamDeRqXDjdpgcBe1odkL7qO+6QQeAkcRb5c1P6x4Fx8QH2SAARM
cIE4BuRKLbCJlTGTtRIuHObXDiKY82hxO0YO7fscBuwKJ2PpPF88XMat867RRZDsHe6QsQ+uorX5
V8boqXWm00bTbLdq28QkpRUWrITNvnpuMiNBUPMA+Aa9bWG/9X5sz3Zhp6kM+o0OZRzLgTrT2ol+
QE7R/mlWAXvRI2Y/NfU8W9G5iwzAT88r+ujzQYx5Rf07dqH8dIsljUGiBjEFdzNzqmFpftdsHvqP
cgdeBw0BRNrHGSfwGDe7oOrtOfavxyty/MgjzakvBx/O1UWLKCbTl1fHAlG5U4p1FgHwjpwObcSM
LyFrDtT0E1IZuLQCkNSmleYWvghzaY69Lc6xa9Ot9kbFSv2EIjj4Jfflqd/StbKsDYh3YuL90po2
J8injpBippYJMQ/9LXYhT1XRAmf+lL9DURfvdOc+0mTTm99jpWHeG86sFW1YPQ2+yJUCUYd+/dZx
1XFfp1Vt5b6PrvkbUS/fyDHNBP2IwZsNi9Dkm1duPkyRoGMUah8pNGbwKjcnK7fmTTU+1pvcMF0a
P8QFkuyPhHq6i8zVl/o3y+MSPC1Lu2dwfHsnrfywoGKKgNLBx8UGZZ6KzZIzknhUDqgV9MU1Wcr5
w9Kdp4gh1cvkG8dNaji+e2YTf6LujGnr7oy6PWBmZVFvNnS6O0m0V9UyScLXdb4ZWCgLr2MQOboS
3JahztNBlsJk2J/8jVnIhIfNLweuXk9ZOOJiNgeKLvmMmPzBGd2BnJ68ZdnPNPpNTqgkLruKw/Oq
vxDqzeAwp6VJiz/SwL67KoykHbs4SU6tTFk2RgZoO3gqTqhvlcTi/B36OcYYrx2tnD7eluEHhbLf
AEmGRbCqrmBU7ZaCBmjMupR0/ULMo3e3lQd73N6HCrE3o1BawS1WRSHl64Fw76N0RWlmAwkurcyy
grBEjBH5OsQZNkGqj0Dk6xTbjIK7RJ9fDGT1DmgqlmR6RYtou9LtY3Y6rOeZF7ESdiyx4TJoICYx
lfcqTSM3/azVi2Xl+p8zhCj43pxJd0BCMHsp0SKRT+Epe6ct8KMuezy8wZOtrLvDdEzGdfPPQEXf
sGrR+AHBh5uHhUSQs4MGYKnfF7Lz8PgchjYwfD3DXHoPcwlalMqkU9rXvrq4+Fx9XO5dgW4ww3YY
mvitjHPoN2gfVKh4Y2iszvpc75MMaNcGgMw9ZNws8e0m5o3yUYlN+3aCnm0TpV1ZQ0l3bqCmH0m1
Xz8D16xOr14Kw0InUHT+ppk9/nOox/RY0GoG8Sgh6P+poetF8oqiyRh/GlBNzNwj2cF2rOJmLS5i
dk5eP/vgq3/DYV7jyftpe9NDXXZrOaF3eSU4HEgZb6mEqdMNRFPoSxA2l6l6f34UnXfiN7hWKDV0
iU47sC2UyMLU75uB9Du1G7I/AOttGEJ+YYYtS8e0tR8AF4OhYI5mr4wpFU4J1JonEC0b6g2dP+if
E8EP8lEoGxgwwPFJ+u3EVqiv84AzF18N26H2+RoPBFVrOCe5QRkfHXFikrvSoYlajx4yw/g7+H2X
9b4U9Npa7XToghpd+/AB7txFg++E/WmLf+muzLnbs9AZDPfE4pq/Sfylh2oXy4dT2uuCetLtfW9x
tq68plBMCzeVJjcGjXXQRTifTxkR5hC72vGwVUMQtXv5F8JICch1hZT/MdQvSdsBdhAGvmfQNYRR
Z4AjRBE3e6hfiZPQDAJb6ln52dsCLAedh16d48iPLdc5Gb51lt9gog/75b1RNPDRottuoFc7oKOH
Prv9p49vX+4WKGL7EATLpEFTG6hN39jBuMHx+LUIYLulexkepe1xqQ4e2hhrOJQudXZRv86Mu3tG
aRenDu7vdY0zSCjPJ5MONFTVLXTpU2MkuY4juDLJRDNPd9IG2kH7FAEwrp5B5gYd6sGndttrjAIC
MHvwzfW9RtAHa2F3WxPXAhzi2IbTwYr0UBxJsp8KdW6HPUZL2QA3c0Dr7HRPEqP8BJE6uqKFosx4
N+XMax9OV52CxMfUCcO74tQjOD3vKnr7oRIT9GA1LY6NeTDmVaU2g6qVtyEgqeEIr8Mm7AyyrnU5
Cfv9DFxNSYHBhtPZdy7Dz1z97/06bxeFe5524zv6c6xsbk9Wfr8PsfOu1V+wDwbHkxBQ7iDcwl/M
1ppp2sjGcSAk6hGDRUTB+4pfmNo/CYJHR71XhWuK5cxp8A4b1Zgf33g5PyUO6RGTD79zbn8LDPXk
sir/+zrR9gb7DnbzEwe/sL6BhbIWbyIsJE3LVWYxK9C+YcgIzLdfg3At/1L/oAnQ1obeU/tRXu2O
V5aUzwVH7Ndt1KHhKVE9S53t3AMry58jFiMvA7BoWsYSTaw8nFecpDV+i2XMicvLFNVf3DcaeFzB
/8J02Sy2nVyD8ONI+Yk+FdJhr37J0BN6CEOxlO/mvhQ6t3cBDBsnFGvpBexpDsH6j+hiPPjOIQSJ
KT5z+BaH+w93PAum7Tq0osCTnf1QGLX8P8EBv55BTNsdlv1owJFJrX/6RoB+EY2+kug4YxhjoSYb
FpBU0si2UD5mpRrnLa1T7GTE0ejY2fLPFdO1i2oNvOWg/f9v02NAXjxzPS4/bx1xu3zze/9CgYsc
2DROnw8/DSRKHT8ANmAb3Q2oN6ahof0EXWqT5LbGMqRnLlrPP3xwmQjKVpcEBoVX7r3xLLqncr/u
vz1zGy6AsOtzrIcWuY+ysnBXc3+k1bxOWO9kfwZoJ+viAht4zJYm3AxrC3wqbrrqxFnrPaO5AeNM
vKa0clpiqVae2CtS9nZ5aVWuaf1qjeDxphnlBXR+um/A/W6ypVKcbvgCanCJ9o5XDGKX2Eb6Qnoi
82GpFJ629MWMSQdOFvaa0upwLzez8LMXogKVcVkA7iB7sUypnLlaqOwlfl8WQ+gnH3SMdJIV5Gwi
Anti6p5g84mO7OkfHlXrZE1kirmB1KIcWYONhUgyUyMa8+ZvPp1iagDo/DwRCjc+pPsPCI8Sd9tx
lMYzMnfQPBePH77RFd03YOlK0FrredRuBYiFKJ3Gea9PM16joPea6QHI+2Msd6ez1SweSc+9IEie
G9f9WS4RPmD56AHg9Ev4rIuhxWT8PVDXrFlhTGoNaVzKVgrYbfMl9KvshDWs51BviCMib6QetzSq
kyqPUH555I0AMqGziE956TqhezWaoUeP+WAbkAgr6g+keiGtBLt7oYMJL0aACtw7vMNi9qvZ5B4x
NLwrWu0c1agyfv6XdJgQYLNrxpo1XjFLO5MMQv4YLGbzG8g79CkrMu2FUhviM+nbNvnxCTx0cpQz
dsveE+t9hTnNWCu7ZAjUqS+G5z2Btg0CwleXJUqZSyzIzE3JebN5CaluUkqMeqLGIxlZ0ZAFzyHg
mQi2RTtje+d7/skXInnDSnnK6x6pRIBsE+JxN91r6jRxsVN7hSNWqTPHad/lEw1bujb3rboUo1SO
IfMXZg5rHwBFRX2zLS93fUSoadCIxslJ3erzJm23eJ/qPDWMs34VtsA6e4hiROe6u0Q/jjp11QGT
NM4H1C/mxEzXsAifpOXIDUK/ZkNLIVkoXSDc2Y5uf0VhHebixm0UioBjm6jSNitei61IFBYXOK/5
qFm4MAtyqKcWniS3AAt+g7DQ21jnmCBHKuoL/BlkSOxE6LNddu5QiVNjzZ/rSK3a2fUsqQCyC0uK
L8tOqBKNBZX3etqLnqkOcR2o1KYOP6oTIdyG+uydew39sGHtL/5mKlA3S9nVD/vTAOjbQvEcvMud
RJESi23Jd0VNVjY11mwH+wFzNmxJGZUD6DHImg/0GZ8AcBtIg5TBAk/ppaCnk6x0gD5ZRosubffq
OyGOrDOWKYqTi8RGmSuioYmcsxodDlRnCFmq+WygAtSGbaCbpj1BLNxgSRINxjXIFr1Xtxtbb8QB
an4zZP2Y+Vd76q+Lb/gpncxxEH84WNrSxBBzpYn7p1YkdAT6w/V3Qhr/aGj1a5ByObsNZEe0l4mN
e8sQXtSRQv9dVNsjUOCWhIBg8WC2cVPFFj7QXjkUQX94zJPmC9+DRCZg28iZdY/7mcrizAb106ha
7L7mTYpFG9JacTEOjgRDHuF44VfFn/nQClQt5p93UIrd1hMiumVTaNQ+RMEeErF9locDeWpIBhB6
V2caQRVL9mqQ+wYtOcOnzG4THeoYVoThiOVuRk1lz80HWnTNGATkzHjegFc1LGd0yYrpdSUbOiRr
WunTsMCQyPnPyK2Zw/DMIkhGZb4sB6+tpgLiF6y1+OujigzYIkuJrvda6ifB0YQYy30jy/etc32M
k4mfCTaHWIhImdmjiZZW4kJBDGXwybmQuC+XdQbaGWunDZvhSmbmFHlKeGlDTWBYiRgfHoxLIzf+
U/917mHcCyP8yINmBF8CJeXFWfG2iwpcoyLNMV/OECjzoAZHMdB08OiKx5gKJSm6W/fOaIHMZNGu
1DFa9Tnr9kv//XRbz/vT/GoQmmchVhBY5ketzlIZzoSIejsuy/l9UXjnj7XQQCC2G9SyH8EUJnO9
5bjqb4f9pcPsbRsfjbAeRpfyJtDW0AIFqAzFGRF31ap9D/CYDo0apDNvexrAPpvTmfsAUoohIkwY
JY32m0z0AJKOHdK0SnXChYhgik6yQEJ/KGq7ge4dVMqWhjC8eQQetPUeyYCPVX55HMxBFtV/EMap
vesC5AqVoxY1LeelZmHLKhPoILbFZmxeR5D0wBKZpE1lpvcVynnEWbV+IBUHWFc3nIr5/EypAH8j
uk94BrQ4C1dqxF+07WlP/2qFVkNtu+hUFOFNwZf+oX4O556ZhTGJJn3/zUWmM85J+I6x+AaXuX5g
Bv8A3DoE+UHYFCkWRxa3JM/47H3LXGx4Wx08NxfvjsqxaItqE64x82Rvule17X1CJYE7tS3Vr0e9
ZFOe1XjF0v4uaIodFUhyocGcOWDF2JW1nJa9vwdy1Lvg2Ja7PSt8OSZgXU148paL3EXjg2/zUZRo
d/oJYZLS5NCu80gR7ININgnrzFQAA1qDLHhvXS0nkJUVFx9Ruf4W0KgJDv9Lwx0bZydMjruxybRV
sgNDXYbf6mX1ougdnfA05YSmJ4Djad26Vjp4sSlgID+ozoB7ROOUU+riSpeTjJJ0cY1SzByV4N6C
KYGVexWQTNsBx34UJMwrIYBwtytqqCjUCAgS8qkcZEOh3fgUbl2F7zIqJ08qgYzX2b+NhJCEHWdR
ZcyA7aktFxSC45xbfjYk78ktljYuQ+4fHvdb6NS+lHR1ZApyIVdjoBjZLgBeZDrr1GwL4iwt5MaE
1/GvvSeltqkWii6zWp9mk7VxsuCv9wdiAHRFx/takhuwR2T4mHIQNePmmcAByX+wzRQQ3IhYaRqM
AEh6iaDF/IJRbR9Ss1BO4L6O/GyzZ1AAdmY70MUaMcgpttjKWankuIBXdp4ryctnECPU+E5wtGuL
/MXgizukgDPgUWsE9hICmYKRYvIVtklj4A+PvxKNhp/ejW9mqHNVKDWWF3yyCwH7xHZZEgNrLmey
CQgdhqX7LY9arkkhbvygm6jsNuv/QBhrDZeWtyPHLFD/vUGA9dUWLh04chpt6cc0H6/TuKmBacaX
h+VCIDu/15ronuSDOSCr1FA8rlxRAu/ZpI8no+GJImNZVzoj6r6ApdHnjLcfwmvUtbwJvG4NHiPz
qoJ1thr6ntaoHkpRepXYQmT8pp3RFlrWMF1WalXpZ4LEUs1vDl3rLtDyF+6wnNb4uud+CK9ak2OB
pHkkJtnq8wvOHvk3St9v8kg2Y9KlvRb5bIQZGlRmjymPJmZni3IqkfY05osm9RpRIfw0A0ogkNEf
GlJtFQxd4Bo+gA4H4Xv/6SkkJcL6PMwyP7NYuYpGIM1+24H9MBrA6hfnZ1M6cD1I2/S1ff3HOA+r
FYjy6wr7ZWO7CYWokCDUd0vgLFMG/HeSHfLtwe/6Hy3eTXiG8ZNyBMGpoCaNGZ6WGKNKe+okJP/x
VXNZcH9uVmNx0PBGD1f+8PD/PpmU5J6HZ56lAwwCs6kjXXkEbrLe6tnJBP2zaadqqR6IlgxfudTc
4o4ecq0zDMxlSRuxef4QcsSwDQpYWtB5pK7bhwOs5iPDNXQ1cUuQk0lyMqK9ylk4ze+NsEon45Dx
wFhpnXDceTKX71OPdEXXxrBwQBOQZ0UuLZaUYC8YSE4lokfEck9fkBiWRsdVj0v2DshkhMBuR54o
pnH26ibzrCHWD++9Tpe+CP1a9HvYAR+YsKEoVU481IUYPON8QxMhNexJZsjXhpCzCET9vGLX8tzn
htEAqG2gk6riHpLE18JMmZnKhN9yPT8g1cfOK1TOxaj/9/uFHTeCWJQzsxylVQ4znC0Xgad+Lw28
U5D09XdvpUlpropBQrH1U6BVuMMw/JWvcNASJF78VnbdjBxDqLgcE1areBJ94BY9Q0THDYqYoxOF
TTYoYgQ+ysW0CRIAoS8RPx4qMXctwG8hAngsbsRYhhXAIlTk6y5nk58lV2dbiYUwMRfvGjD0N5zX
1IIOHnJ6aqAkGxWV3zkYhP6qUKDV/P2N5shiuqFkDmXauBJOeQ5oBoTaqVtbtaBLl0W1HZsBa5XP
Y+lMoaNjGtIHiPY5TYyqfuwlhxDTn3gZokwp03pU/CmxAc3l3bRuLk1XMlJoQl2qfU4LVvYnMwG7
97wil5689LVpIXmgCbSPcedZmiLkyah3DutFfmhVnpChJ5QxaVoCbJkSf3+vTs6VGN5CPVtcsYOL
fMDPdsfAsmxGmK8EBku5fCwFeO9BA8WlAgrLmUM1jTbIWOmz6Z9olESkx3B7OV1BcnAgL5Ym6pVo
9zriJWXesm5z0jD+7gtWqLl1wsbFq0Y3pOpVomgD5ekk83316fe3wY382KiVweiMIqFzfjteWcE7
sGBHLemymcqiZ2T5xLxF90RF6hcmvon58lUULgC8D6EIBJoXrAFYH1As2Ko3E1LsiN7iMKgHKSKT
2V7C+xyHND+ED42+c0rDRMKz1Hq3Bs6JdkF1dHAfNi7lf+WQzwl9LI/aSCmAHLkO14qoRDSzjGon
+nK60BRwNj8m/CYZO2SFD596MiMQeKsL7dafIEmJxmntg5MzsRFPVMRi61j5fZY72nNoxJuNU2AT
X6TdoLMifBaAXKbZxlIRR8mz5CuTdgrDjGBLEs4O98bXY7NcZ7HwBe7Z8ldvFQpt1uR6GutjPZEn
Mj4A10lAhT6r7aKS4WlP5hxD7+UpeQjw3AOToswcW7czd77kT3+HOmR17VqkNJg5LU6UmW022aUc
WtLPYVAVQrhvCupCKEl8TRUzjXauLx/er8JgCV89iWUArVcNXhaKikdKlaHfzawEn+D3Tj9U3s2Z
6C6C9oyaYn39VqjgRkQr/dtVcxBPyIUFU48FmEPHHhNDk0+z1cV+ZdnmXyRu5tKc9K1pJLRME6Db
jdj7r9Rzg6373Q+Ojr+siW/y/T0T3f5CyoJUwBZhMWZQP6r2XwbGP36H1ZOZYi8zp5m9yi7rWaPJ
rabgLfSP/P5+6ukS28QRUY+knOtMi0uVtOnOFWQtQ5H/Vv0A7dLsEPMgNp+C1L93KGx7wvK9UQB4
fp3gDr8QN0oM9VsHNRPYjM+Byk/hV9hiAFZFt+59zm7s1gTobfZkUhQGvkrsFqCheFE6kz0CrnRN
M8SaDsQ5T23YM20/aR6FxM17vuZoHKpDrH3B+xVk/jk7dh9dKOBppEkR8LVNeHjfujZuTc4ihPms
kwLspAkgz0lPI6FDTYc/7bXQdcSiAA9vVxGTmz9oCI+ZcWfPwLcevZVAGhTLXtzoo/bE7JD9lhsX
TfMUYZxYIDtFCoFcJt4QpHCc3MlOPrREmszj1DKhNvR5kTmCqpsPXjuR0UbbmbJmCFcm8cKUN0iV
ESggl/O3KDfTrTk/DwkQf8vT0TXbkWYLRWysTb1yumSk7169ACrYXRqi++C+WHnFkGWFVsxS63kS
394Tzu9A9f/QHkNgrF3ebTnYYVEFfRLb62VCAbyqK7JXJvubsYHnHGmfE0qmA1n4ruJTaX7pRmmT
5wDAZct+jjb+B8I4/IV0Ce6M9HIe/bF+qWEsc9Kxpi3kHolwiNxk5aMlSFFVZm386Xm4GCsWc03X
qYQl66dUH10hu7ySr0MWZrIx8/5L+YRXFYBxisVb0RxyWdZ1+7oRqDZJNsL5hVcyXyxZK/1J6p0p
HBMGw3Ng4FwgHwwFdZJ9laSCtivSqRIVubEcqofx6yyG47pLhlt0zehyu9ndDNhDH3Sb0CHF3dOd
tc1tDsv2sr7rx4cuQZ3NAfqTa4hs6v3qTmRXDJhT1BWbfYDSgj9GsmpHjtgdpQ3F/TtRs9y7vyYR
/BSMj89GzaWfuV9X5SYOvsi8/O5YtJVNQje7dS6yRuTQzdRtXgEimbTkctXFaujMJ0M+nOuxqisU
iFjdX4IAtzG1rL+zkUdfPx+UrtO+CNtIhwrwEjxHE3a2A8ymf2IGenstyc9TZUKPQ1/8Vl0L0f+s
c0iF038XpYX9uRuA5SGwJlj4dhD+pQ5RxuzFyzE98sLraE53aNkpNLOdLVrqMw1z4/aUQP/o1Hpu
1CJaPo0kke1cD0ZOCL3jPQeGLjAIniaG/pjveSuDHTHS/WV1EtZZETpwpasV07M064D10n1XXQAW
m41JJBzpZeRCi//2cRGbuZU2gUZVh3Fc/3FKtAX2zJxrmi2gEZNaCK6kXwj08gT4PNAL/3Ukqjkd
frmhnUOPnv3+mfLAyUlTWUKaWFE8WcrQ1AWetTIth4+OreKPCuXe9oazm7m1fZzmwdMkPwTJVSE+
DEwLKPpP29EBbcI1f7pRL4+tT5+wCGFusJz4wE5QNvpfYwnkeLRisTriqkyvakbzzCBim5Z0nDzD
pl2T18WEpkEaioZKUliYme/adqNMQiBJPKJ7Vhs8shTPr4ebp0kb8KDo8KV4hlsDFMJldBDPt10O
VbA2y9/6KHAvgk1712HUn2KbqYBVwhu45sqJJ6Cxe7UpU5Oe8nGDJMlgx0uUo1wgeoyhyQZvundV
t7LlAuWuWLn1V6vzQhucI4Xc7v6Zhf2VQ/SeKd1rXpfFD+i/Y4XkFHnyS1gWz0wFDzV9zy6L9lKv
YH9B5DAUHEtDrVjo4Wp9g350i/zvRy2Ne+Kv9ndxMXAcfR8PCRCzrxxJ9wLdLHk99z2/9jjrHN2n
2YKUQSOMY9+58NtzJnt41Q+6z3ker/0/YMJaTwCBQV+D1hGsa3NgfVIlMolh/pyzzv8u4ywU1290
BUkchVetJVX0/KQv75OjdkPqOkdIsgggrUbNIMoPKkWQne5vxrw7e6M2eunRyE2kT/fsLHsYVXco
Ot0l25NL957lmDKaIL/qofuDOkYdYp+njSj6uDRV9tLhevvKQWRfQq8i+N0fNH+x/Smz3G8473ps
XPRSwPMT8lKqEkamZowf41UsmbG54kHLSoBCz0GbJdsTm2a8URzsuWRB26ZXPWXfUoEa+gjyDPg0
rUmmYgABEZU7sdWcGg99rcPzBGXxSvXAyg40v2WHoh2WzB9TiNVdPwtPcwwyE1odBIgOOgRo/EzI
CYGAymGfvdJFPwFIyFOVQN8aJDM15i3aM86kIl2Py2VlQgz/0EN88S779xwA9lLzor3MQMkrMwNl
wwQKAeS13X4SskipFv0CIgcw3XqQRNEUSzhTaQ3G/eWf2x9rlY1I1HxeKyLpxBRNNZsPwy6rPmAC
iYEo9RVpjuKsJRn+EpcXz/ysEuVr4BzS32p8GbHuxvQFVqklu7CDa0+xGb2gwqpTCGZPKvOAmNxb
SpRo1dAGoxa4dm5yHNUzAcf4Y9mvyat0ioEA56zD0ykogsqI9Zyf3UtZdAhSPsxG0UKy7fit7Q3z
6DMp4CEyZm1d8GFsFe6Db4r2esE9AeCRp9Q0qk6L/3psmpaDKkahE+xibwmFqEminniK8KDfFiNQ
CgqVn4UJOkDJLEfOfN0nphiEGAYfYq/RV8ITJPCiiCGCnjumkvoz2J7Kb+M3TxL1VdcDaOc5WVaW
aDV/vVIHx4Bl9t1PQ9GA1Tt+8YkPdHhNQ7hvuAy5Wyb/dElBhss11xQu4m17ZjtE0VYSreAGvwFw
A+96IOjLNqn4TnQ81N2WYHYbYEZ6haWIxCsGkSe/i21gcRg51OYJ/fPvOqrPbH4DW3NaqiBFDoKR
0ROO3YMZYmqbaKyzaZXmr5GQl9U7R5GekVasq5Nr35YXD1VYhpdeSoC15kpvnqlfqLOp2tPCJ1d8
moYO71Y3t6B6xkxjB71iiAWgSYAq1+dsney7Dz1dcaK9ytmJ9E4WShz68zqBMeZ4G17yRzJF6TIA
pra3DmK8JK8UFJ+g0zSoJDUMc6OVny6jk0hjZFetF8t6EEfcZc+HLSxHo5uitc85CNZVPJLeS4Hh
D9iN0JRg7YrVTve5mmumyG9Z8bhGGzNPptpv/ZPBTKLjmbLRO/CA3vyUsRcJ6znSLwfKDNMyUSak
yrVy0ntWTQIDStur92huBuMQOWjO92SRR002U1Uk9JyS2WwU9PvXc+42Znbiesi4U2AkwsDJwdMm
CzmHVf/828/QRs/c6TFVsTwT6DPD53DO2MTeD0BbT1nKLy9YXmj52Dr/R5IN06/QJGSTg0jk6pj/
+96MozxzQ1b7KsQ4UXm63FNJX1VjNVrVo/gGEClsIABQ4fppUW4yGzo2yOiM1ouHvRriRSUhCTta
+oQ5rJdJqoyP/DCM/AxXS6uRj0wN10oYwFu8usYwL3M7Ran2Xjr4PiLK5VZyVg5cWma1OAgwFYz+
k/Gxny3pLkHoBImQup+sl4qXm84DPyzGdUo/AXsuma/80vY3IS33MtYrloEra2+c361DlDLNrfr5
S01D6NGkXz5xU4x9S1vjQedcC06qVkTApDgiUMTSzYwPKPOCA5iOrxMzz/dgmDrQWNBxiPfIsAqN
r1BFbLzJqOtCkBJsfk5GdBc68+IRLSZGhs77QaMld20cl5G2Prwz4QvYkZ/U41/WVKxfVVWOn46y
Uf/7iz9rgVp+/NqFs/nN2BAgZPl2a9uLaYnZChn4BnaFRpvxeUwwB4K7EHu/fAXPzZBAAvPI9fyz
c80rA4aZTk6GKfZKJrKgf+5JR1o5CX4zlLGjv5fZlQsOjhOdwOG/WF3ltxLpmv8KWhBNx4tvzOEW
mqkbW/Iif2QFoekrFlvuIX2CO+ITUOnEDGsMe2ba2KYGDDITP0qmksHdWGU59cUKj51SMkBlSJ1+
iNTaAn6mqC2d21sedcZ5QG9P0HbKzxQimrtufO2PJ2rpR4m1m/I6DzIQQ+5R0M72lW6hw1juPCrE
DLF7hXE9Ztr4fQdp9CFQSEVYGlwnFVS1JnKiiHNT41LMQS2IQMyMjgzhXxhj6Z/C/R2cJed6vGZu
0Cw4SIyPv3/bccWY84jN1u5zM/oHMiWXCCiSkbxSMHAqV4dIJB49IqPi7+UyY7BQGPrW4owaedfa
AYQKcyP7AjVs9teklwJFfecZ4YgbAGFuR7UPbeCcFm/MfuK3rJQExk5kxsK1E0ndtxOtkvXyKCzG
0Afwq6Kdc+Deg4z7bfKUOjnFxc5M7h3VketeHkR+Ag48FRgeBc6wxCTks4/TUbKIIV+RCrqmOkCC
AZPFBPA3mDCZkc+HAIz4kv8MN0SONwIV3DB3W/3Xtm9UNwIE1R5kE5rlRLKzFqoT4xxFuFqw4/jb
2SwPO7t6Jo855mR9Dq7GJMvsVjBVgKrkd1grglaraa10Za3yjlM77dhsNReYSmX1o0CKI9HM3jsL
WkclUdwUy4uSo1asqcN9VvE6pXokn0dunYFMnZtOJQpJfgoDvGZjAIIxLBbWyTH7tdn5/76b2ZgC
Y6BrW/fdM4wvqF+MwO38mFIOJ63KoZREFRGRjVoUz4ngY1TkaEkulGbR/pivcQs8haPxCLl+L6nv
oKjipIJ4brsMCf/+AkrM4Tw50DUEcPYdQ6YyTPvg+W0PByTFEcGHqanTAuzRzx/OufLNO8ttDEpc
2kcqB9JCnAjTIJrG3Bb2RugZalX3PsaqaH4va3eRTYPTMoCSncFNKt0/sspSEwVSAkBLwBQqpgRc
ts1fDOvdYG2JWsakTq+02Iq3K6bHNWJTJ8ZUAnR2cT+65yHdZP0kt694EKG8GutOq8fLqQjFd3A2
N8l27MbSaEfcX+CR/kRPfhWRysU2fT4XvTXk7spGTe9M3v6k1g8EUajE0yLlpxT/vQBlKzrWSh/O
iOgpG5p9QhBZacYuQYahMsycZ9xibBN4jn3n6SoTy1Fihxi2wMKECZZwGRu1jQ57FrQFAqPk+Oel
RNmJRwOM7PDfh4acKNmb2lFOgygUMls9ma9P5yXJcEnE7SNahA2BJ0VmH/zmZZ86W7LJHjyHdIO5
6r5OBVo5ak7sWjYh3FybBhXqbVshnGoXxU64ojcePFObjpw7HnLs88wX6Az9nBvadWAxKVaxu7cO
uKP8kHYKHEu2WS9uT5YGWTuzEm+WONiv0qKXFXetDDzQWURfeMWv52Wu7NO2eVndeBWflXk0NARV
VAwjdE/89xSzCbA8MuywJc0mJpO2LDTgf/e7/Mf03YEGZSu+mp58jt/4z1PUwMBep72Xvjt5eljW
fLL00kJi7/nSebGysRs4QAIc33/YNPiWlpLq9rSUNUrgqASM3LhZ98zsuvSx7O+AzzxyZPIQRNB6
shNtvv6xtVJgNI7YWUho2Wpe2jm+gC/D89eiO/DTZzYPr+l9/Dt7cWNT2JRxglBtNlP+bS1n+TU1
NtHMgl6M3Ch4QkMBykNaQwrUYmnXmHsd+NG4eAxax392CGIrRmscVJRZwvoeJAkUBa0013s5X5CS
aktYA74ZVxNUQA8DVIlqOx4v3q47ohYwP7lTXqnbxiyodRnvlOpx/Y7t6/eZYP0699VauZ2OzdrZ
Jpapovu5kQr3sQnUG/3Q5cgsoWK1kSakmF9do/Kggqm19k8MI+IJ/QaXzt0rR0aFmo+ger2gLe8H
NCJwyoMqIMoiMeVGRnSLPDrqJmPfBoNrou0qIHKd7V78ecDVrJbRNrB7YGxsKwxe3A9B/aaAjFn+
9LOiseMqjPBQBuAKFZC59FF++LqoL4khuvKcL4FhOpdU9noG12U0hWoqcJsC+1kZQLH0GSKKmT9a
TAull+uEanX0YsDiKDpK8KDmHUDxivokJhloHm16EcrcUoiI0pJIHsFdJF4K7iUfaCVfZtORp6Uv
MsDfCPBoCKN0FE9sAATX2nYHOKiZUQsFZT9wEVDnhB7Wjwy8OYdnYUGiR/A3E9+kIwrBzREe4mSE
RXOGvdFdL7wxe/6W+yFWgkYNr4v3priQgIfNuQ/sgAIGxPr/cmU8DqQqYElxFnCTLTQOXiHpWbRT
wF7OZ3egcYwYCRZDr8Oi3XFpmBQkyMI7RpbUkYX3kSs7qRSVzQw7/CNraPeDv9fd5nmFeW1T615w
yo5wTmco23oVNOThb2U5kEExDaCLjK7P6zlA/IioAOqfmVE+mUc3Idn5WxM37rmzq8dsh0OoCCxV
gchXYp3XLo17zT/U2Eecx4lMVK/agafeLVssa7Gc3ELwtG/zSbu3B9CZW2ubBhvMfPUPdOIjPH+s
Ons66Kd8Zwz4BVrYNXYodwz7y74eJYg37a+uakIRILxF8fhIcGtVO8c9qEWgASMDLDnTE/yyy4FR
J8Z200y/hhHvVnIIo0jYg9VCy+NZ0mAsmxovXrUshOj7s8SDHdyvJbmOwp+hVQQMZHMOyJmJ5oX+
QyXcraFqlawsrtUCL5nwWg/5CyehoAkpf+KSU0AmApu5LP3Q1Q1fxKWhCXF5vQ5wxGT9xae3R6C9
B84o80Irq7Fqy3/SGY9V3MQjjXeLvu98sLFmlP2FxaC8rJ2yAXG8mnkeOEFOqvxguqmDVzMOvSRa
rzckxB5Q8ejdgN7aEhE7GiEx+LtfHp3XLI5wLfBEZqcAQMA9GtGqzb2QU9WGNQ0L7lmIWGd3v0ZP
4l85Wf2+YKnSo2tsnYKrppJ2CSiM6xxzK1xmrYur9rIX6/XEeP4IXsP0uQl7JjmBu83RScN8KztL
ABBvGQK0J/2pOOb12MkKqnrh4OuOc42/GHhaWf5bJaREUlmK/7E11I5JlgT3aLaZCc19Hi8nCP49
OW5xcNUnUEj+wpquj1rKpr/GAuQaad1w2SeZzCGJZDGlGr+12sTxTTN5quNpBp29xqOjc/z0xj7g
aSaYfKzE6gwqPGKRlmiPQ9kGhcxIl99t2l7qrg9svgc7HN8mur/6yxxZxd1ShvrvD2QfyAlkQ5xE
+v4OssLNd6lUfyPTKnOOnhfUaIpAyGz+UXJQUJjI9jLnvavz2XIG/xwN9X0zEvJbYk+Gw5mdIuQ1
wjB5rE4Lwf/eDrT386NSJkXLQQy+IKz+Fd8fmS9yUigyHzQaYGUvMRUBKmIJFFSnie6pE46lEDLO
oeGBgRqI2ABkEUpK0VA2QLQ4yDSdvRx/JUr/79Y+1Mz8hAS7EEtj7hl+uhzrsCaAwYBGhsJ8y0e+
vm6mgYQUiy0Lsg3uPuxmbCot417mVcdaeUgoAwRzrfIPcz6EJ+F/lYysiy+DEWdK2zDjz8YEphuW
Nin4re1P+/KoLyAYh721WVjU8wDg/FRafTAUdGVxQnEkHEJnXFQTUoLCbA05cIdU67U7CBMc5Qxh
EVn2CMtPhARzuY46bIFZPI00LX7aSAeoqLa2+W92aA9l27QI2DqzSpfHO7PDSjRs6jvzvyqyKoEK
xp0a6SE1x5FF2UIPxCeDq+P8WzZe8ZUS8YOkY3JEekcTgZzVur0teLd79QlH1gRizMCw3LeTg8CO
K4R0G6H4m7a6AS3BawG6wLrSEAITuHMJLADgQKTIPT7m/8jrzlccN/H1fSAMN2PfYQ6NFNFCGolr
593gZYR1v+hjfUiKzCFi1SOgn4Fr6fjSLns8liW6ObBKY4m/H2frE9ftsUc16qr1R8j4oS5/krXE
bS33bm8j47VcC+FwAzILDJZ2KBo+jV8mKLy1ccDujOxZ2s496pih9nvOpMRzQCtcRmZORI6YvkFE
932gxhaIPJzD3UbO+K6oNxvOQOY6nxkZX7kZzbze5hrypaG+OZwyx73HVrB8Txq7Xb7GdQoQvfga
KS53x8KOy6At2UBHIy73G23n3n3PjO5shyEU77nr7gkb1QpmikfqXBzjv/9nfjSCsSMd24HiY6Cs
3oabokU1dzyh8yplDBEapYEJ+RnKfj7pATVXth2nCgvYELQZs08bsYcJCD4AfUQRHwmkOjEBTs6j
h4eu61qKx8kCdo75f9de8uDtmxsLdLt7HVKjg44yobLh4Jx142apH+zw7ZTLcHddP6OACe2V1pE0
oLddNcqz1Z3vfLQuh4LokTymcGtTKMLQbnJ34CEhS2lo0L6z9RFk0ejdUSH2wfV2g9rDMsr6fsGf
ZhVNES0ebWfrrRmr9yuvGGC1k9pshaSPNWeKWR4ca0QqZNM4sqs1cifawYu2N0U/DGBlNTfN2396
mSdUjNIx8GTTZaicr9IztbbY+e6H31CXuP4Ab+A6tQGKD7EWWQk8y+b0lQf7OmfeBFNB5tNYaPKi
UU1yVyOjIO7vHaagm4+rPIOBP7caV15maHDmgopfWqhQMvNESaQvVPkYJ3ml8NAvaNhSjWWLQANo
gORB0mg9XraHGDVybG9KIOFn8Zp+hgOQbn2UzpokiOMJxtrpKGE83+0JqvozpaTSHsPytxAmKaoo
yV+VL9TUR8K5wG+G6Qr2D9QUwkU3qJrxfr20GGPL44jnJ4DkAcOzMc9NC5Me6lxhaWOpaDoFiQ3f
h6WIaVm0r6DD/lArdDDRMMh17aj7G8MfoD+sHqUDvlak3+HkmdkvaEfb6uQdcDivRYlYh4CEv1E2
W2apLFYIbalbXm/CAVurV9NDzgSyD89mlTDc9+39P2M/HKXtFqarrB56pjB4G+QtV2iQ6jad04A9
j/Ru34tY7cMCxgF88szu10a+pAu3ph67p/HTctJZYF4XI8oDVSH7PHOB4vhHehe+mxbQEDxLDR33
F8LxxWhzAmFqX2HbbW1WXj27r6Y2T5G131p6b3HmsKUzvwsv4oNO94QzrtEkP3FUXbtENOKVS965
leZ07bx+9/hINkyLqoShI+OdT+RLoAGyzLjL3NdgjmMzFBIqtGc+ya6vsDW02h+vPheEzwjjDCWZ
troBu/Y6SjBG3U+RdzhdEmmrDDtxGWWb0ulqWGAuoBBtpOVkG0jS7myXb07SWuNSVNM6C+n6ehUK
jQ4891kmlj42dG3yc3lXFnKQ4pr8TQ6exo3tXbW0wEtPskWdlDAxnWpVlMFGfjL1Q/Aob7KboUEx
d9kA5UHFCc4Ju6szvn2g6SY3DioHBMxn4LaKJX40jBCOR8hiscyW0HzCqAPs312iSkE5lERm0bra
p+K69qqhD2SKIwWNx+KzVN6tqvz1HLsr9+xZ1e2X2z07ajvrRmIBCrxqBQegupfqYbNFonGH/Rml
Q0y4kvBGKsBxcwARsGe8P3ppGUt1DeCO3bQBrQFeoKgsyQFlaoIJP9xMul/9oZYlwmgGUYy6cXO2
6ms5/u4Hdo5ueY5E2MQtw21mpZUREqxzJrpGrSU8TEV1f9ElNPsRuRulOTAq+BgMczpwwMVf/HTG
7KXU68So2J7IHo1wl+BBT9KFtO4u/RO/CK5Fn8o8cskHSiNcZ8VxToJpcF5/OrQnjOuPIsybdliR
ygB0QBSkbUm8abP13G2hcQzkzRN0vruOXqNQCPJuFo9TP4mikaWOlVuAlgnFSN/iTWUkviFGEDx8
oJrUJK0Iw+j/tVHyBl+nn4bOP/z0zpROJXZE7LF+f/n8nmg7/DrW4oOFVmqJW7j7KeLl9pTH9rPd
jMP0REzjszuLYAWpy+7RGQqSUwUmY4MRdNoxlZPattbLirBJFihVVLz50fr+1hs5nQ3M3RC41vbH
FU/LRXG1F93g0/+UBLQgYsrpHi/76aJZ1GMmqgrNXywZYeM6xOeTCsX4nB/okloYblIhDzh5PZWc
kg02yahmC5iZprQPEOGUwvttyPVM92iRNhFoa3qZylpT6nGhDFNIDkdYmP3ZF6LKrv+2DZsXBKdi
HMEoYiead0I2e3XEQovG0oMA2PmC48FF5pmKs5AbewaUdRgLkqH0iLYmIoWpgSKOSyks/cC+4YLJ
QCL+7cNA5Y9ecGC0d5idUfy5y87WLQf2nwjhSFYnMLdXtnKdOc4+41ucoTk7EWCYxgB9oFFpYMEK
h3rOMjZAhmnTXXLazxppd297v256rHrZpURk4vVZJuRtqlY0QM9RNi+7kBFDJ52LPtQXklRZ0ltP
kOlS5zZS2bg5ihLZJCFS9aGbDMrWNo1my19xw/gCRVlaPW2TUzmublJFX65c94o01fD55ksNm5/j
ZUl/1fYZdEwce/p2I8eswxezxpVaDRWPPFS57GIPMVZmivUrz5lWdPOhp7u1HE/h1SuMbmp1OBjB
q/nxQHvtavbCy9u/xUAGnXme9TnbUZR35a+eJNTjH8LfboIN4vsitiNKH05lCUsuD93Raw4CsAFN
HEsygBZ3KVrLM2801sdW6UZhGuzCGt7lLaqDgJquD4ujWEMp7S11yWah68rUzaAxmJiMC54HKhDS
H8oi17swx7vkm/oXY76kPUm9c8AmCjhbAjtjwOZqdrqcrwRIE6iOqUP0svOSXbMqq6xY0QVGFVLn
ZSZY+v/cMkgdYNneHd7MACRSyEkhMyvqNWWW/ouPXoi1D38v+BtL01ekLzVR7Sdry/5hLzNGJuvA
qIWKZy1p2HEri9Q8a14tYvonERi3O+N93O8R6wlvJxEPZ97w5r6myywyYJG3bDMO9Djih62KG3h/
tCnKgclmzjN+nN3EogH0VSvXjx39o39pVT2aEFEzMGWM9LTxPk84QYG6N1HgnuAphcfLSoo08TOp
6Ilu+QM3JUIozBILoYuuVEypar5+ZP6k0MTxQCp781oWXFasfUDSXvdgCijWkEs+wfBYEEURVuY5
0y0wILmk4ddM7Jw9BhtodN6J5WU4r9sNctA4vy2qHV5G+jGhZ01tzR8OIvvtVKNUd1MGddPOm/7f
B53C6W99jJvmzVrPqK/2j4v19lD35SOB8cxY72vC+dq/FeERvGZ55gX7Ojs7jzJvnhr3tYbduZm4
GmrCojLrZOAf3SjArK5PFVEMq81F4lEC1REaUDXc2cZT/VmkBdt72qBAfAqACO8jaAXpSxtddSKv
AaDUFIAJ9hRhtxx0ub9K3NyvV6yrPq4F55pvYkmuIzCgVjqiakxbf0Db+WSHN6NHNJISPyCTDuKZ
qrESxIEFkZQ9ceoY0dNuayZ3msWYL6gT4zbhywpvRcgWjTziANfZrhgF8f8Q+4Rmj5S3aX+uCL52
Ao8/O4TTCX5vVHpkitYmmw70cdj6qZOnSFPk1d0yOVqMqMNzc1eBfki2sf/L7toalWqIyxD652f8
s9RRFqwzpHIsJxD1J4I9/6f4B2Hcg3oDHv5kBs4wjmAPnYxSZH49D8FXni6BEI8ZhkIEYd/YfUBT
2QNZ6BdpD5RVR7b+/TZtn9ZQ9t8CZPzWXIrioVUymNdmrBYY4dvQyupDKqBWAmUaziOtZeQCKh5+
ciHgwtlzG2jBc4FG0JcvhpQj+Xer7yeuH5UMLuGblC9yJDjvbl6ucqfvgIQltDXJGPr2ZWZf41n/
RQNObhn2eiWwmix+wUCZYRNU03eDWTZX/QSTtV+Tm0kJA4jLR4ffSSl8jnlKE8VteKWddtgwO0+8
80QxPOIKI964bEbskTvt2KK/rDL8QjO6v+QKSZqlSlGar+wTJxmspjpFUFuWNRLuP05n3xh8auDG
goa7FmzoJz0BweeFlgLt8LZXCxlcdaHLqnMIKvg+RJbRLsODlAgKspUE2+8ByEIlCciAGzZHNoFL
K7/+scHCqTnXIwA6sUY+TarvBnak2tJ0dwrS38DulvJMXobKVhAc+5eFj7cGJuQOIt1yQRBZ/1zC
WuSbGsnrPceIry0xbISTUgPKw746DZD6rlCXA1022S1aJOasEtqq/4A7Tfy7TBrPRqVd4PDwsJY1
RLX5W10zskjIPwDaSQlXetR0Zo7xVYPkGfW3mnahTwuCQW1xnP2J0s9jbiBk5h1WL150TJ3ymhF6
r769IHIOJOFa2o0t32FkKCcCKv/efCSIiU5ZjEcXBoELeoU9tgdK9uYGhuYfeSB5sho11M7H7d+Z
JT6tnZbnBEolxjcDHyLexStDAr10eP+qNTHZYg6BS4Tofpyn+URfk2kdFKZ6Ttul8NpwnjVD+R7R
lUBWn2mY27nRop1JFMghKejF2z08kvcD7vrioy/eHSX0DV6HxEUOi6T0YOtCFPZZ0zIvgzLxUFp+
lF2MvBfRWaeX5BFbWZX6WsUhWxsWaXiGhRD3pVtRIRWgZ7wwTxPSC0j/hQ8gEBDElvRlG1xmIhBX
SczUj/q0xDIiLZl2wwRabw/NPQ+nYEplYMVSokqOqZbj5pYdEk4kZg8VAV7BlM/c5pccDa6m1msv
jn+OtE6V8DDEcl4MsIcC8cQPhVsu88GLUYBtSohCue7nV7YzvFZU/sB9p7FDlvUMv/MqAazeh1PI
Ge3sDgOCANvqkzRb94+U+m7v0utJn56RVDq/mdQnc7AIK7sPMiKTJbZi2/axNZJ7YQ1KvUqz+gWw
NYyl/8pi9FZcIPzR5Yk7gp6CO5cifCC1Zv2U+DM4OThHQvOzymPV+TBCrrbO1TWKlPU5UGFX/6iy
9yRMUhk08Mkzg8jgMxb1b0W3PeeRmyw7KQATIXeeXzM1w41h9rzxRHoMHUs3RT+rbtkVCGH3dAUi
iw08RXhTF+Fw3VxkMdg3B7miqjwJlVW47yp9STEpiXqz24u5YILAXqCsjw5WQLnolj7uPjvaDji6
yPLSpoxgtFzp2BqYe2zs7l/QfnWAS5cRQc1DWiTEW31Qt7L9/9/nK8X3+mEeWzPmB5S6d4WeugOw
mY3quW24Z/LHtCwvBLz1GScOAQabSTIT/Gtqnig1AYoOEuM3XCN4KCPSpPeMDAmSPksczWNO5ao0
T7Ndnt1wVEHsf0Prq1XLrTQ+eqAtPfzPVd7++ciDBN43UG4E8cm7gvVNPnqdMUcbK4nDguoYjuoe
KF+Iyht2E7dnf7garkRoulrxXhTrqCWWiTVTXkjycuxyNjUXYF2pTwR6/zOOgZkEnTe5eBz6eEET
7eFCnQsN6Ob1qjVSLqy4Pbv2OBLjHEQa54EfiSv6GUqoHOEcEpsd4OwBj4mokwelbquqSEguHvhg
r4yy7V8eu3chsLfwDFWe8Jl9QQHlJWyQFNFy+3VIoT/E4bvCd6Api8DNOr/kXsIeH1xM/bXkxumS
O/Qb7QlR3to2FGnmoTjPxAQ3ALXtWMbvWXJh2eqMKzCgZyj9Dnj9u1amyw62OzqIhDb6obYU/Ovp
cnrhCLLThF+AiTjq8IBFybD4JHIwfWuDHR+5bvzax2jSHD5r4FG75w/jSBNzfHbz7unnx2vAqDEo
pkhZb2Y0locCiN2FnYm3FJfCBJV8tvLLy7cbnUAT08VQWq2dJmSVylCJHziYkLRRXmtyPnU0n9aU
luwD3ToVV1KafNlA1tOCadotuEYEHVr97oDIixXpCvibT6K5UcrJ8Dv81nE2Nn/lxBcpbXCjQO+J
N4zqkpdSTnwAi2BhAw5RiRFTf6oMV7IwxNCGtzkwC5RgLfOj9/ga4jQ1Ju2KJhPUyEPlrbSk8ft5
isym2vjQT+eTgL+uY123XxV3F1DXsiSpu9by5M6meHVUGTjbLLgPBidKA1uJ7zg6bdYJAvyuZOGr
GO4bF07F+CM/KqNo2fGM4nhViC2rsYVJAZ7p9/8rEWeEfgRedgqzbfqkTrjrXOZTuWKPQ/zN6t6D
jsYmhUmz/MvRm7h6881F4GkM1e6St5ZdmLkp2zhoNypnhPg4jUb2MLPCewA/edfhQuQsBv7Dchbn
0y0fzq6gcHrJWLBGaTZxvpwOEjD+HPU8h5EpLyH6myaZqN2yJUJEKfocSO4m04TbmhzL+TSsWSXA
pGyOEDiPJ44r1OaVv/lLPhG2lKoOKF0Yx1++zRMvDYgaMzp0J61cnIfU7WIrO6wew9MmzATt+yo4
HaWmEt5riCLUY55/zs6QoQ9TpMfrWdRGhOT7lDxSY9BsXJoYfspGG5hwJqNS9f6dVyR/+iXeH+PD
/cdTegDueQPQ7r97YwFeBUSIlH9+P6xnF1sGPsdrFSyJE+7fc/3PLtYT3GxiEG84TmMZoZzZtVY7
6ONDpVDEDQic6O5YJzRc6H3O0Mg5chAUeNTqkRncjv814mXBtzLAOvffzvVg5048aARQP/jQp/Up
talHkmfJri2seWswbfOGUQbkNccJZ80XrsEvuxkoFgqIkktUJzqA+gwTPD8ILhQL9jttfm1Wv0Fr
Td1JmEfP7q5lqaZxEYlCvEeX5xflXdpKygza4tJ8p11X2MWtPUHibnNmMNO04xiVYwRN4GSFU8tg
h6m+l16dFw4ooFTXFimVFrD4R5Y/pFDXCSqxw3GapZEjyGL94thpr72LREovlfUK7PtJO3+KWpqS
mjf1CgmgKoU/AdpMiX2mZLJC7b7X3rbjafQkfEOtVLJ/6ADkdxPwUeRRz8mAKXGh+6qeAbkjo9dH
62/bMHhByU1TMK7kGRezwJ5JNJOEtdaZXL8/4TUtKkjRJ/XO53h1jZKdR2CSbGHxpT/7DsBhALUf
hVZMlnrTGtqzTdtOz4MSMAwJL1It2T72GpMfYtCg826HXE+fYn/5+Cuhpm3KEVbRakv10K79jD/F
8E/5RwJWhu1bZPfvk+6l7KO5rCkTySJ3aAx2IBEahQcnNC/GKiKJg9a2tJSIQ7Fmh+qLwQy8wzDv
hR3vb/90BEk0ntHMG+NzdNQ1xfSmQRUP65Z7JovkkkcRygJQ4TFuHEoH4gkNshdfEO2XWl4Q47AW
wC5sPj5EECMx4mHboCBXinRmgWNnZx7eYLwRR43SaH0DeHQeo6xKHgZHdbFETUV51XDrNHkIp+pv
OaK4Ae44P0eA8AmBc9C1I6BvONbw8aSLISF7LQhm21KJL9reRJ6gh6NuoTe4dAwo44pvuzJe1Wwy
JHjV2dRCcJCfHwFPmQB8GP2yCb8HS3HWj4E9xT/YLCl0/UswF5DJ8JTJooNKHaIeAzX8T88zW3ew
EwkHm7eKBtl08ymWP6wsD+HTM7NtytfXYcgw8k3NM1xmrtA+85KyrO1zhXaDtdim98Z2/bLYGFT5
Vnh6VI7cVoi+YVlVATUi9BJvjYQIVz27sYxh7JAtTFRS7EHa9ERXd619wFbmarJYeeChdae3Q6Gr
1/d3K+NRJKmD6r5JygcXqs5lw5Jpv7C11SAlee7zcaNpqYvpVmnG60+bdN05lTVzlSSQhtBuvuZO
jDso8SqDOMmspsZBKRavTxT2vO9pKPpsG9IhhULonjbj0WyrIbRDL1gEiN8nDvVSkKdy/h9ZQ1Cj
Z/yM19xQN3NxhfI8sW0R+Gr26VWiQ89DCQTvd2kJbpnI6bFnryYJ9Txq32JB/AKjbImJ4u9Kis9n
S8IWDmkScCsocVR+Wwm6ruZj2+N3LRTXoHTR/Mhp/lPhmiP1cwHMlPXAUV4/KMz6CEwnB6VX+uus
CCt/gIgGPB2Wz7Y6LLxMXS9wo7qdI4ldJHs3YSg8LpkFCSMQIHXeXpBTeFNv8SwPSrqEiC0Ail85
qwsoYLr59EE/nDHkwkOXLTSBhPkNoOShI3gbFpYv9bdnWX8CaqAWzSmbQxEPsv0qEutcI13MjG8J
8TVVolcTZydVlQ9h9sxcQ332yqQS63effySeQY6SrIGBYrh3NHujC0NcjMpEmI28T9H2FpDOiqk0
NijCeXyjVqRgw2+xrBjfkMi0iDbsUuYqGB/M5HjN66FyiPOeJYgr5sJSdPOCl+ko4xBCzTd8EVMi
QPB9aS/lsG02RsN/6Nm9hTPTqjClJ9CtQEyNQz5R4tWv8+3niYCaIvtqqU/KMOIB54VuwfxakyM9
EhxEMaedxAKdFOE0OXtCFS4d+dNVgR/hjdwvtmt/kOY5JB5WyB6jqxvzvkd0P2+Pu4GWuSoTzGab
mk3Ic/Zs2s77IUUoZfs/L5BQlSHip8pGPd1xagHSYx/fwW3oHgIxtCKzxZDNWl0SqTXqsoylXyul
p9YwoGpuZa+otXKZQpBuHlLfgM0Glc23Q3PMNlE1QDUa7loGfvH0i7yMiCs/VHopUiq0BeV8zbBx
0E5nPSHI1QjNyvA+uKgyU4SHIe1/CheSpaT8XG5zvgYWIuynCauTnRGZFheySoPpgl/IpYX1Lg+w
TJuytK7T21J0b8SKN8WHHgH8H6tiCL/+aC4GP8xYdLjmZOg7JRF4TePeY39+ztF9YwDwfre8rOEW
Z26SYKUSqbuObh5pFShqFaem1PfHbhjB4aeQ+wwFke95PaZIt/O4yCO1xwV5a4xTqRlMqn0ewu7a
NrOiElJ7e5Z8NlXQjkyFyEh+qiAjV5vsBA4uo2uZl7G+doy3Drrk0zeuNx76kuauEVe7t2KXHXUm
slIq52kOs6UoFecnDBLpU2KRjjZZvxSUbO2E+/ImAwzGdTxw8PPAQDhyqgIG//qKzBl/KZUX4CJ/
2ormdDMnQsVdGvsJtER4RFMX1npdtkNEkssIbsZ3RW8ONZmDoztLhu04mYKpJa7e3SA+fV6L0v69
GmLSf8oiqhHbtqCOYWpsN/eZJSepnP0q+tKeSER1Xibq8A+h8HADeb738Ad4c44OND1FfntbV+8F
SKJiTqFr3JxV4i6ax5RU8Xbfm5HykdyMv/X7lsC0SEtDWSg8wHOPHl64CZkU3pn1fIeedJGzZvyZ
fwxmkuX9syyj3j8cmuvP+v3ZBIKhC44jFjcchwvgq2Vayt85avNg2wvmlMIonW2YDDXghTtlxj2K
T5a38cCqNM1sHYIJ8/4BGi/daJRFrWoLhgOMROZOXN8skXMZnBtGdjO/ni87Fjv1UgsxXjgpAmH6
OHJp22EDWCU82x4CRXqo0upzSe3/y4HtpCmiMSJh7Kbnx/8os8Y89MKDA7NLQ2oMNtaFCv5tsKO7
Ral6icOPAPdQVFRN5ipWo09MPfLUg6J/hL8XXOzj7xeAdrKYhmrBR4LjnU2pEAPHOSnx2dxtf+jw
EQ5hw1gjHDasb4zUqmnwiIEgZd8EAOM3MGLP5b4SVGBCRcKj4xcug2AD4Kr/5p0tBp9i24CQaCWA
P14BPrB19o05g7WkZrBwX8LW5DjOlzl9fen7qYxwZGJMecWxfdSGDUqEE0yuoI7ns5Oaj2agF+Pd
P91GjQKQnxBv1Thn1OgTXcrpXfHfSctkyxCKney4kao20DtteKg8bTfxN3iFJSPX+ZirnBi6GyWZ
/65lwMQOyBxH3mmOMnL0Af2ItFaAYcP+Srxwjk6HKOJUjfS2OXcYCqt7yEQuH0aGrtkRe81yt9XZ
t1vhlkKbBtGBFXU8Oppu0ay/5GjmXbm1nPO6SMEfRP/chuivOJRl5TRl9dxuC2wI467vAMGogjTv
rUoZcFWp4LMBWrsIBeh3Lxvxy+bSvn5qM4Bb7+ZJ43uz/I5WBmcX6ZS8hnFkx5O9y5ZK4GR2R3BH
te0SEZun/XhXyOOBykMtPiJZgI0e3NtidXjSjqzVEzAelHeOJa4vSEHa9gfMG0rJTR6snJ6+AW5v
g7InLer8BDWsN/wo/HBSM2W2PenLnMH5wYzBVh/OyMSeUxhG/mpBtgMYgi3+hsmqM784etMiCmX0
rZXg94MAsfEmotIUocW48Z/+F68Kh4tg9JSA45mpztbdsCxMIlf/O5unJjHlKnD09icfG0ez/5ky
FjRNt0C60mT1WOcb4fnzzvwkW3jekO0kQthTfOiawX9Ap9SAW0TmBzc/f04pa2hF9UFw++ZdkR19
iGhml6VimjBDlz/QJzWhYzztMW6Ldf88preKZZyTVWxXcLUa3/RNEtzkA6J9HpDHxOJFmr3T0ylD
CJFEB/FnrCRmBXGqBSQzkHKXnYZTgSjQ/0Qm5ckRFYGcDxu9tB6Qn51k0hskw+J9UFVmMHStB/Ct
a5rJk0S/8o/GQucrp088LxVmbJ2BgSl7VLES7LOTUWTiE8WHuMIjr+ArnbBVzeGj3w6aSF5BoPmB
Zqe0Gn/K1uOXR1MBujT/yGJISY43FkDMcVJz8R49+WdpF2emEL+KxPd3jiRhf+N62xegNiEaUWFk
RxFHm5vP6pcRR7pkZWldJpSdUB8Mc0UjFjkDy6aXpsGjoGHPwUyAHBth50VG22k/CwbeV6ja7tmG
794ukq+F2vNyO7uUandJnQLBfLWRL6TtMeQHLgIIG8bP7EabtJu6Vezj5SPx0hepSOd1qqfvU1ov
x+VcCdyLsedRc9nkIh0FfqkXiZEG9FPa0s1ABlSJlIhWXX1U9MaZnxBYPuBtfP/PK2EjQYhtZcK+
HHV+/bMsIuoq2YuaRfnKZGVZSLoaLZdu3m2fQ12f25iKmp3XtxsJJA8HwbzxhE2rV3B7KbKkrTIb
t7MI8wHGMQYBkjGcYI10NcQZRFy6X8TvbojNxDi+eu5Vopabw9ezfmqpiF0dUcYdKV+86uj4SiOQ
ADtifP3Cublb8cSacWFCz1N76BAFVHinY+MDDNJe1IKkLbHilG1S2IW3GZCfSWe3ybUB3DkWEoN1
zR7vfKXd7m57KQ0i7O/L6fmU5Xyp4IgVgcndX5X0iXVTG37K4ZiMWjvrVfTlgl3yNFcNLDNE70hV
Fu1KI4IhpgzKr4UPMQWJjAQDV2jfJyyvfjZvCNGaUfwoIECZSq+ZSXMoeLCGz5yh4YgACtdNYHGp
1O4wjjdXkm2RkVa5ucKMv8Yx2x9wqINShqL/6YImlhDaP+bJZ7dozZ9uqcqXG3XxUBUa8KXsqdpq
jOW2hwkm9kd5jVdxtSz8fF71N5t3NVvT8Jmko4UMFMEBYdCUqFhU4sQWH1D5rvcYWbwsYdaBZSzY
3ooDjJ/jfnz402ZcaRT3SSVwBRqN+tLjJrYtOreS6Rm5aubHeSEnH+r7lD7MdfyByTDL0hYOMaUy
ESYbF8tBLLk2dQo9Ck07rJvv696dD6WNo2gwCyj2+amTEsqKKY1ZB3KpDv7qOJrf7Brd5YjjF9c9
eg2GfU11nPY8J9XuAAoYciBQ1W8T0NB8UBaJHv0TkbbSLqPfpAQ2dkoVr+rqVi3AxnOtlMP0Tifv
jCxIXk1FKqeLpkY7Yrhnq+GXj4oLcnjCj+ZXZVVt9FW9d2IUPwiTC7svuKqlFvqB1GQnCPK0BYMu
3nmOeXI7zP5/8SsAxtLRaPhAgtToTFNfe7KyAtmWzdhDkhN+umnbgWkLnngfbW2TrM81dIyJoiBg
YzVcg97QlaH39MtClE+dvycyrgA1TZJjtXfqwHTgojWair996G8x42gmNsWy+lUdasIte9s7qQjb
rq98S2sp1YTQyHdmK7wf3xL4Scnk1oBbpCtM93TVq+H4hsdfs+kQ7ESLZgPtVE7u5HRaMPKGXprt
f9HXjLzNOnFjbqWtLceV06pRSu0iwr/0brUEjLu+B3xjNmNnF6ZYYFO1+MaZ95S6DhEFIY6tqm/D
PwYwtgf1IKyvtSgWpbo/bDnHO4QOUDlxLHGsXu7ttSHKINwPKU4LQiKGQGSa6koKeMT0f+TNKbkm
Qxu1S3ab3sCM+Chqj+X8Xy9Hqu+cg5S5MoWhJqTrYDqegtkb9l6AaGtOvFxaYmCuikSBUjccmtgv
71Rxv4nIOIEowaLQdaUqFj+ZN27AgqFPuCStGYsIrAy0QO0LLeTWmcv3pi0RR+lbnGnsb8vGq0VZ
pD1izdvmGJ+YKyeFDpByLDvCfLXPmszpnjmIsfmsQpffHpsgieXpjj971EeHP2mmyEabe/2bIRzR
zFN7qdqgSmOh9/esUgUioAN8HlRtxfL3SiRi8rInMZm6TwPf58Ki9YuL9kvZwh0+Bf2p0NuuJc/i
LXkKGr60MRmss1zI87SSXRI0tEFIRa21gaRu/k57dEWNPo6qeUIdG3df+v398GNH3X5TRNkElNbN
gP0EkHZ+y8thcgbJ1PmSuTqwQo8nqmjk9JxwxrDOyS8BubjrSwgWjRodGsXLIP9PC+CcpaR+DRI4
x3Oqxf+QnND++zrCujHHgmUbyX+JKapyVq1YSaDWXguCb2x8bSILRac2IyjffC3e2wNqtzG4/8zD
CJ7aGWD3LVPqA1mp3J8VZBlEZ9QjAYlq8ab7veodOMbdCBgJMl7Wfys9200bjsBm99uJtr3tn6O4
47zhZtiK7Gg8wvSfnox54R372oJPvkNLVh1aHvR6P1CCI6SaCwNb/7FFN5s5i86RTDEx2cIjEnyO
rFc2Fw4ZCzHFuZtj6HQL5TtVorfFp0XmT4RkieNqdteIhGNmr3W/8h6pU1kPFz4mJAH7MyA+vhCY
SXTdGOtcae4ODNQYvJrXzK5CmQHzzMwkxlKU6CSMxv53R1aAAvcMBRxNAE8S1N6fkis4gTRmJKNh
OUAsbP7KX0iNFsyn/ipPJXFLyJ7MiuJkrsO/yh6sWXaB1AnrJFIT8tVnB3P79mYqP0PYm9yTn9SS
OCXw8yrHdxJ10YpcMoi74mpIIgEUY1Ld7xUHpl3kSQd+BrWk/6CsGHR9eBk/1XN/8K/heLeu2atj
Mubu0fI3vpa4NSYmrnhxLm6ac9sEsZrH7adFRgTBXAYqFTHl3tL5ZbtNSeWgEp+BooSd6R13AW1X
rhpJElxEzWdy3PbrWNL7XuZQJxvIUGs2BrCNPkpYi7vlWeH/lrTFbvjhzr9/kYV8GWaMl4rE/DFD
GY84hXPS0/h1iUmQXlKsH2sU7AiZ6+YFbHVC2d5YoUw0JQA3JcJQELZMiKsmz/tZpML49V0j9Biy
qXojuCPq5exlQtrV4A2UOri+9bvW7pv9m3BnZolzCHIYu1S2qnzqGd6626ymS66gsQYLnlCESRBO
oZRM8pkyMsUHWy1juilLU/2irFV1tM6ZfM/30fP/uRN8DrEIq4DnClnnWZGgWVSIGUzirDJjG+kT
RgG+CF/+LEfZg9H302SIWKQaPBq/alvZXrye0LR7wGVRQWKWjuIxL7EJ5boYPCe16AM2o9Os++jT
xhwtWXI/hlVqxvo8fm5GqDyahOcRrB2rAd1SLuYnWFDdG61XGCuZpm2REnw7Sm7A5wCmI+Mjw+Ra
vueTnczKgLTLFM/XcRHL0Ddqh2eK9I8opTxxF3b51815v9yzkDfdfvmgWAxS3YUgqOzeTBKe5wcv
+Y4xvQTQxiKa89OyND0TsPOQjhmw9NqBx7L1GOGb5is7WfOEYMsFIpnrYdxCtdpKa1ieTVrJy01O
nZNg9tYWro7msR6v8XHZJ3w3YtEjfWr7oKNL88k3xpp6FpLFa3Bunky4xkVyYnh5qPSLRsbeQAjV
yt9tNdTBfZwlNuqeXjmaDVCKSgBzwC6c6qsn1XpCwQpBak6KJZsL+G21Xr/uEwfKqEtg8o+hGCBi
aN2GASWvf5BrpmWdsc+LAYa/QG8sqsGub3QZIiyv2LfvNZ45VpAwbYQ+njcyI1gw+AkOyY0TQfpX
hxye2ekmRnl8FSSIRh1GeLu5h2Hk4HiXIAeh5LwLzNRnWPyHnpwm07lBDKuZAewjY586w8LcigJn
lXte+fxlPidTEf7GPUWk24+N624kE21CMzW85rnBa9H3BjP2HFUDVYlCWf+XG5p2E3bMHpzYFOMd
4zZ98w9Y0RfLv1UPpfVy/bZaSmjZs1nS73A7FkqfE834clfglbbvh6cOfBcc+mkuOhWsL/lWACRc
uVCO1LO7MI20QQTA3VJcsa/CvBvXNgaOTdCJQkaU4sif+pML6w/oP+hM8Hf0CE+QekMvTfuMyQNW
77cPxRtbDW2RKggw3cOy7Rb2xXD15ykrEoh3WAcydv34xsM7ujMdM51SBncxpy0bejUqKCW6Jx6E
S5gZTZNbAF5xMkmPcZ6zWANF5/IzgT4ZKPHgYBwaoBi5qjSzcMpjy/EERighyAMPUYV2Qt0K5MfW
aj2xqQSOwImSax2C4w4OvXGH6DRb/U2GqAPDMjhq1G5VBN/Ui6O8pbtMqujvs2ICaEPYkLcDhmqS
lGr6V/kTrbSO3WosLzUangQAZiqkIS7zVZbHveYcvd/CdWIqBvsNsph1PWEimzH+F7JQgDEA0jxF
XfcJ+lpIHRpqcBhyizsRHtJLr0m5xtJJ6VkG8EWFXTNppTJx1vg9c/410xlSXX9+f8H+DA3WI8wu
vZ5VpLndZWIu8eEHAKgSJjcyO0TgYV66U8H/3S6B3Hwvjy9K3VY3Oj8vaazq2ePB90j9orjbqmhz
3JrI10DOclNokEbQL4rNt869b2GyPiqg/3YIHXxi4YOslCSdvwSVzyELWBHJDDh5cu76jkdPU7QK
TL2v0FGVzafLxE+n37HUj+Hk28NAdRsMMeXJqVajxciViObQ5QjWj/UZKbuZPkojp476uiFmEeaT
/ttOVmJk+XDQuqDGGHiPKYaO4lm7RfeIKxyYuNaXDtchRpAlj8i0lNYo7/gCmd72jsO0HDCNbrpT
QL9P9z4cBynpcr9rWYxUmTAvQtuSF5UnfTBWTY0J2f1URy3nFOGvDQsCn+QhAk6tX8Cwrx1CMWgi
iHIo0kQPpfouHwvnDd4WTRp3FPlgZj80SjdPgeyoJLOFl2dcKvBNul4FyUt4YUOV9rCRhAzBWrWu
7pAGjabbdagn8tTPE7k0D0hpYckYbwsIkV/8gb7cnPkb9zYcLTrf17/cRbdoh+NhWi1OucSTnxCO
pnleMc30S9eJiQEVZ8ck6jNyFtvgRnis/qD3UxgW43SbzrL1r3jXirlR7HVx8JemAHo9ziKPRIbe
kunlsHgAviYrtmgtirsDq62h0z3XQJ2JHBf6tFcn0mvh6t+GMgYHKMsyYpU/4cDLOgXTAfsqSXDv
kg6JqFBGKzXYzSmrANvEfzImNde6q5oLWKS089bN7aMUnn7AXambmpWuRpVkvkUc8+G0URG4X8rs
yNXou9m5OxshuJ53RhSQ+JEzGAKkvMRYJEbNdQGalleCHMC3Z0pxysbfnpIr40Xw2RerVb8n4GSI
gxIrT0/LicQTdErDfQI2wfhHTUqs6tH8xSEag6SbGqcrrRlM592Mm0nRQXnMHHDs37oHVzNxfjNA
zWJtwMbjCuejgVzm1S6ri6Cxv6McRuMcLnTWPj+FS5TiFRwj6A6jv+f1cxOM+TBQ8wglQppzB7az
fcBgRAMypU1rcPkaUJ3KQd6hZWGumJB2k4sJ9Cl/XIGs2bgJTK8VZPea5QyvnrJ94DWRXQtqhtE9
cNWOJrxG0CVN3LO15N1wuGGKyWFncBZqMRKa+DroPR0q7AN2//oSFROh9pdIhX+Dmh6Ze5zmDT9L
XYBP/uQKJsgJ48ThXOXveC9cs0Lwccu8vs3HU6Cp2DLOsWYqt7O1rlBeGAChTrv4HMBf+kf0eM2g
oNvLihzsYVrssD03l0vfNJZBZxpvF/hPnVpibk3o7Y7/qO35Gq0gUgE1UG2Bd/tLv1vbKpn0VG1j
STwnI6bTBEUVSkmHdcqMMOEk0BxXhU+3p80gfKi/mY6mtjmnygTVA03hdu5ElfejXWhOfnDjSpl6
DMfwQY4x0WtbteTGv+wHC6tvXFZEOzsPWlvDWIGQ7NFct0f1FrsBjg1M2TWrpxO2zrPPeggb1PUF
OdkitldskessJl/aPKZa4XQimQ4xcNFBwBlKG33zMT34y1J9MzOsKZkZpqANCEWdor+zCTprUfxO
zRXFEQh/Y+u0B1mk3yimMycSn6Ny3wz4b4HAqaeJawYkRkTgsAutNxKqIjphiCQxLcL33rMybAF0
efVG2fmFxs2V/1U6F3ByabaXUXypoy1VyXWoMDwfPvZbJnn9jEOgL39Mane6yM4P/JOu/CWPo71h
pGeee0nemvREddfuTugXvl1qdOeJRVLLnMut2SebBP1JBNz4i+LC6uLSzQCjwWg7e1I9qTCbsSUL
jkZHX63Dg/FZSiX6xVFe7v5A8VNyYDLUNU3O9W79krT/d7p/qBStKH6yiWDMRjKL6r19ZwgTcjZX
QeAI1EwiKH8e9XdSmngHcE6PNyFU7Prj1+6KqYOgOGj7hMRNSw6+/m+aHPDR/AeAjyKtt+xbcOKx
kgBvXjhrSf2eZYIohNkNJBw9Gv+z9QFUBNRj1oWiSM8ftw/rwNQXXbMqZR/ZYPA9Tn+hbsHuU5wb
g/fK/BkHwCzKsYbKfk4Jhv6zk4rhuM4JCtAf8Wy+ppDJqNukzMyohMbKQFUIF7DeurHiU6Ii7PT4
knQcmXE/deXerOoIgSJdDXQHlYNKO0Zu2dyamOuiSxdbT9Wz6ianhhvaDvV9eFIrJbAkSFX9Oqcy
Loky2cnpFQ/1nVI5QUrPX+cDlvuH9bVYoZ5+jwl47kMWjBjR7xc7khwU+4zvE8CvM7dSs7Vq7FB+
YUYagaF2TWT64w4ibOuDwbwV3XtFL5Z2OVZlpA1jr09xnvuhifjFDiT//hTX+AfxaaQp0R7qsl99
ItiinQ4GFXyJKbdNoaU8vvf128APmKg2/UtYPOy41lIXuWbvA6fAAuCnFWWnTQLDSIPpHtY0pDdD
66Da+OKbjy9xwyUEqhqU8ysr8jw9Ur6AC5uDDuMfAA7zS32BM+DO0yXGntUze6J8uA/JNS2pkLWf
30wM0HFTvqpzWNH3Bh4bt3kXQo8pna4WkT+RO53fn5Xb0DIRlxPVvXabT0b7kUTj0V3QyjpLcU7q
PbioXOKjUO/PkTMnB5GvIQoFq5ICtMD4KdxneBBOUzOysUkN+pRxnBNe8fO0WyHqpY9C8et6wecP
6e4xICeVSjFK+ELns2RG8IIP0M0vbh4dT7dmfh/0F3nEK5n7lDB7MdxSTf0bCSPQp5fKb35z5zmu
KxAK0I+QYUiXc0QEMFgSQvctArkPAQXQBvAD4jijHYRe/9dcJNZS2S+Rw68wdDRbHxk1Dd1LBeyt
/YTfb4L4q3is3bL1JbHDAvooTL35g2EwMEj+5l5K6K5ReBfi0/PGihNliYtqWnrrzXN4Z1rhO783
gdcuI9JhqtlQFLHZlt7GjuEN9rMdezJ8M+qFS8FRl35w8yLl90dDCyFTEphc4+cMRT3jtBXtIXYV
EY4whR32MBHnhcdF2CB7eD+NykMkVzCUTBJTFvvuVV4lWlOh3TQ2CJJIXKMFItRFH5HBXQ4QYGL7
U3vTprHO4PHrpdROI59LUxbqXwLhnyNp6baeOIth8JrQutO32SMJ2pzuprR7z6l6z/Wiw/uKOMly
M0Ho7PQeOuEM0Qx2lnEcu8w8bwfvhtWDp8NU2py6Znaamnttyjk2GcD2rmOjq/LeQ2fLmwJX3RD6
Q67VpDBsNRjWyPF1KiqJazVycTAwcpq0Gmdt7UvNaQ4fFA+LnrAfsAd3wMPJ9vJGVmuw60mdtHbu
Fjotu64Ew8PSokPBnFsIPctX34cFh2bkoAfpolsIXSYly9OhvvOjHfDnaSPm6E0y/QY6bl0eMzWz
hbkOwMWumApZRo5xPis0VfS7eYHkism+xPD5XL+N6QLFrLTlqJQKJxlOnzCS28pS9uy2yPz9bPtA
UgqZSIQq2bYUd5xlYggKh38Bmh+xl5Dg0yKB6Jp+n3Hv0mw31xnFnEL8RlmhXPMTJfTtfK4EJo/W
Gn5re/4dO3KAm/u5XEe6KGNV00PtvGen+xZequs11dkbpUClz4rlaPTOjN7/h9megD6hZFEQj1cw
msHEBGuXjPZa4JXXsl0iOR7H9R0SP2GzEtQnE4d4LAIYaeymlscVc+e5zrveg1h/UzTErWrLsG5L
z5KFNKWDoA2FSFly9BIQsJiM0RBWU5+4bg/xceU3sUeowXEm7b9lMBfg1/UdjTdWyfUkvj/8Am3j
VbUjWeTBVONL0IOh4vJjL84qZfuKGYeaekknbI4rBAaeJ7PT/C+j65AdL1r3r/rk8IHofaWJau/x
lounEk1fCAuEZmE01GEC2xh1xorpbUFJgbBvsGRLcfgm/6l6UWRRm00APRgjJdS6NZVdkW5Oq6zX
6rFHo0V2tG8TH9nlXsUS+DpqqvzVoL37pywb002NOaMLjuKAZFPt4rLrIctIl/uBs0ZwibKj7y1f
VV2k1TfdqzD0I4LcYZUVG07+0i4JkDLjnljhji1VoTcn+3uv8lPNJIVqXooVqS8nvY/oId22vvga
hBeTSoe1YcgrAC9UsZpy9Cdi319NJCXUCQKTybCilvf7OZOLGKUVPKI9tZiHAJuJoihNDTLGtjgc
YEj9lQcmKuV8MtfltImauwS7CbRaFZaW5oIwfTiPa6Ct1MbdJjd138x6KoFiGzdVxUxvjavHJTa2
YZcgwSCcn2UwKgK1WsJB8OHUdGvfvcUtcLP79u1mYxVHgH78LPEoRp8PnF7vL+vmw+6XkLLNRc0q
cumRDNZoECpTdxNrIJw/Jk/X88psSYYLLCuSHfLy8ibbgFNUe9EaPI0cU3xKXWxY+fWo2Ai0YhLH
76zRHxhU802s+r79oRe/RC5TdpbSiyeqKMRe2mPmlETKOs+DZyK6sH1yThrJB4ucPJJ4UyJTn7N1
rneiHpdWPq5O/BuMe27uGMY60ryojycBORllOV30Yvji071uKVcx4gTq4Ek0bjd3222d3q9XS/Tx
2zOJHxiBeQNWOwHKHZCQdpt3qMdT9bT/Fy7V/Y2vR3fYiZrmsAJB8uw4iF/paRCRwd4xEn7jXCi8
VRvrJ2zxXJdVnAKqOOMdTF7nytqadE+uUEXxUwQzDpe0Pko2wOhI3CKZ2xekDObYTJ9+GJVN4nMT
foMhl4UONChKaiNDtp0jJ+txNlEtpLvnKvS/FqiVDgFouN5P8d9N5FTLtOPWuo42VpWJ/0YoFuO/
lIRwO/ff1wp0TSvvi17f9+WYzvmscKopF5lRy1RbI+upKcIyQnwbv5lpY1xEk9N+CQGVynpXKT0E
Jdza3oR8YpgsS0kO8Ussz2qUI0NF3RIHw3swdvvVJuimODiVt0FNXkOwpOmwMle+saTQzySSHzpG
eOUpAl8ZqYkME+7iYVlu7v3STRt/xrpsoqz4Oxg90PG00mjh/gze6N+8NjCm5Il3gfPog40Mx0ke
yL2VFpD3GpK0EqRgIsHdhFkjNpLJuoHVwkfWNdPB9Fpxs3K6GdaEq9lT2APbPJCMGGtLjJQ5lkN/
K2kxNKxwEN+0S5NTf0j7mFVmPWZIEixsJVH/97b52yLzeyOfjvRrIZju4hNkOKyG8wxljI8lLq3+
/Tk+3P4RlGxBcAcHJD0QL2CNIFOiYSbaaF/Z75Cg3WbgzAXGzrVMnNUXSOcbO1XPRv3ZFGKNWoLD
aw1Ok6SX5h6ZGpUgd8vPomYMR6ewf5o5K5ljUbVYOHOjadk4UIhtTLv/adAaxr0e6TH8SkT+cqTi
MSG50/8FNFlFmLFMiMiyfEBvWb/mA1BDyqI5ELKdk3zHeI5KFAnvM8qYMwgtHfjlG3M2TZDGvezF
QQ5eBICkQIFQ3MorM+GPgyfBZCOF6RUMqE2qFNg/st/Ed3ppJlqZW/Wej3s3jsGy6MYOGGTqImp+
qeeBeAfrwcQfnx+BollKNZAaH+3BV61p1hvcMTSOULCvlMIJYBJGDORizXLgTFSLsZ0JfKayg88M
IL+9B623K0g+BDi96Ng0KdNKuMKPBjgCDKfNZIh+0Ei6VY5dgcJ+D8h5xGhwM3jOEL9gp1E6w+qQ
rEGM7xKWpC02DXOW0vfhXYdlq3CKS26ZhlAIbexCIdCxiMhDzRinvjQFEmtKlcmlxMbM5nsfZ9/3
iNi+GzVrDfQH0Hlu1lfXcYi/Ld7Bs4EDg0q3vgL6XlL1UGwwJs6Jk5gOQxGzQ8eeIq+P0Jg9nA5W
ytnBvwNlltdruNnET+wG+mIKtW2ME/FevPxjHuW52ErWnUWTVAAiBbid9ft1m9J3h1ML8c1dvSiQ
rkV59/bTplCYdoh0j20TtNDUCo+2H6sqTJZkzA7P2iXcv4tUG+v/rgmOJsYWExncgoaFcilPBfYB
Vfcrt3PwFNI2j1sBilzCpZkK9VCZWpzYWX78rKAfCAxHNcj6btrVgu6DDLYb4oSBLLg+ghl6Wf8X
zvnDOFll7u6LMr8gjSlSlZLU6qTDd2WeaVbhyTbclWLY2Fld1rAyRwpkJ4vX1lFoP9mmIsfUjrU2
vPiw2FsMLmEGclCa+FFH0WRDaybIp2U0jyJsrxMmQmmmgKMAaW0liziv02klfvGuHvZku8NnLirH
Ros/rhmclLr12vrhrajrrEgPtmTLQS5XMaWEXfsQMr6Oqs9aIMADvs8EmbZh6C57jDjbcoiex3Lg
UF14FeXEC/A3IHU9dJ0doZpD9sL6+El2WMrMtYVvtgAD7g0AbxWjETA1APgO0Z3a01OyxHucC5oN
F3BUuQy9PsPckE8EyRfXjTgbFj2/4FR1w4x4DvrHQfCQ4laG1930TtSHi7Ts7rvZGqloVhV48oRD
Kyfb+sU5B1/HLvTp+xAyjIhFqAi9F6aO+sVfJbiv8PcMWaw30Hp5LL1Yf5pYYZYcDcfCYnQTECZh
segm1Q9dil60bi+5K0tdrRaQKWXx/hldXwPJ56XI4JDijEkYVqXaQZPtONXJLGWkgpW22ofJ3aVv
KbEinwtIkhBAS9hafHk1AG9oAN3S+OSKhMwMeGXdgx4XLTo9IjDBLmnn8cdLvRmTGXN8J8T+iSj7
7F7uOaXOaRFtwz7v7ByLGwEDmIX9DJ5UoNUwflJ1BfUIyq/AsE4NBd+jLK2dg61oUUt3+Qoo/DsN
QWoOySXvbw4Sx9tEhPkUmp7IcOPh9vwJXEAuHdEOPO1y2IEtVXiIG46NE+fPmolfheX5UifPBHTz
4rONyYQBi2F2ZyHMiwIjFXk/E4opLkfz5W/pCKt2zxWa/5pZX/p/Sf8S0xHu5upkJ99VsTOB4zwS
BW74dR1iaF/6JklKC/oTVzaLM6gnskYVQrnOXv/T+fwWbLeSq5JTwbtsjEO89imUPBHBJXCFXUqR
2O3CD4sVcWyBo9WI59NBHABTFpCKEKeL0wlTCWn4iN/hzOqOTNS4Hwi9eFAJubBXKaXeGbpEtB9D
Xqd7491XvqQWrS7moWyl17ce4fgTOLJTQxJDv611ih5Bz1bIfQT/Gjk/hRf8gqEr3HplQvfDAcxq
6dwdoNqPxxI7U7ctUXJRhntQ3Oc+U2zp8PfUDEvbMkZO+aWeegDwG2n0j5Gw560aBgpqPuf6swpb
LiDkG/KPsc2MosruzTH4g4i3KxtJk0l8yZGnbMv4O4N+4sXaOZ4AzoFijVtK6pn/kl5AJuxYVWWY
LMjyNCVvEo58VwT4uTyUHRZiJ8GmYCpxawncIM5PX6hTjmht2wxY0FYqAV3OfHckuDchEYv7jgzS
H0T1pk133iWMd7gguVEztslJyqVFZFheJwnph/RGGFSZEpM4IotYPTOZbSMSuEmVBU5Gxd332hi7
hskAY7TgeDIW9DMqfulZC1RrGk9VMGsjdERXGP7oHBt1iu+OxIsktDy2XrKHsRGR7/fq7jRK/dan
onx9MWm7S6P7b806qddajWuBBGUp6fvNdrz2n2wpaUVjT/z8yYkekffvRImlWunhRxB4pxBROCJ5
RMN6j6Gfo3HLocuDTJ8x58W+Q3cwVUAiFkYgxS6YbjgBbiLZbjk5BB2T4yoH9gCgJsLeMf7TVqjj
uvjBU8S83vIKC88OH8yokD8AS3sKBf+yFhOxVBXSPnL2zN3k7e3XyiJm8atO5TW9wqy0yfSsfV5k
XNGtZn21Qz+PJi/KlIFzbz3SIWpkeGWn3p46LqN/9oxXGBhk5ZhpXBPhwI9AoMLb6ykEZJfuIoAv
aAIXi8quYj1ye4kL7MTPzWyJi6VEdDHiV7dsAciLuZeoInSKUQaRAWxlN+f4V8eM3lL4mhh4xbqj
j86Bnsun2CttBaqLqRUGZhCCstfNzf/qCtakbcuy4xVe0vTnk9qZ2pGtvI2UfU4hCP7/dSmNlHLD
2gr6bJniRwv1GGWTKorgV8YvPwxTD7Rhhry14gNRCoNs/s8i8tvHXQs0139J0BJ4YaSpVFJaaQJ6
jci2OS+DNCnL4wjva/jfhTw1iVvU0jf7ssJn96BwH70J1NvQCjbNqWoa3mg9wmZwMnbMpO1jZPWn
klj/zNL4ZI6/g8BsjOrfi8QHg0k8QkdfKxWrrVgUmtKymibT9CotZS2Mcrn2jJwgBn4jsTrNCieJ
wUCvYT6E4ccHYjevO7GRwJpmwITnGpTLVPgETqKXOmKI9zpScs7/qhWiXtnFIek7fJdc8ubVzv+A
snwuEa8Z9O4CZW/MA/JrVHk/xVDGAD+v0zSyZO9MpS0X8eZmN5MYD0jSmF1M7CL6QIcxPw0wYZ1n
Pniw2GLkoUZ1R6mIfaCVb/H/HMHp4Yw4WKQs5F2BMoUKx2XZHsIDfr5Yt9z9/xRt2DGi2fnDmBco
wct6IZHHC6aSV+UpoNr1XtW67wq7mxGShRk2DhJkoTfX3e0iH/Fuz+mtQ+GwvrpG8fN17v/cpSvK
wwq6nzFN0EFpK6WNO4anMM/c+b3sDxRnF/Gakvy3SmVC+yZhm0KKGttyWAgdQj1yE4M3GoheSxhc
q2+hZ+z7DHH/IPJeRuN02Y/T7NY2ZdW0DVJoY2krOZRBJfWiE+xq1oyjEX46ctTVRjPnWmCMeu3o
qqff2vsi+kQo4P0dWHCIyQluFZ1zAY2H3apRDVyt3NdVlKElNmP+9xm0y9ZYjvAjQngDiD8K3mDU
KQOBxcIgsUhrYZk15bgxpQrsk3pMklN/+bxvj8RAHC08f2MMDcK66yTrxo8Cp5cOfxaMG18zQgQS
43iuSL286PmYs9XaD9wdm7UuC0xQI6IAo4kzGkN4eiN3vHAN39Ylqtd3vqw+YoA5gGmQ/uk/YAfk
8+ySI/BC1HoZtxENJfsmGNmUYPViyCNSOGMaRavXWwB9/Jg/aI/0NJRlE9ZhFDfALQ+1O4ZXgn+n
2rxOeQ/Jq2Eqizs09Rn43MwNpfZZcJmRN4itF8tKLL4B/KUXo6qkRZoEa3SYlDGgcIm9Y1D7DPrH
fwGuHGfvkrXOUfTkM0iN9gp/DSr1DGdgZvjZuuRttDkBRKSwszDZKkmyZuZviU5Jx8/e0mZraJjo
TJVyPw8+mHheI1YPjUebyyUMv6HOXYWAwiS73WkVXHtBzt2zhVl8NseNaWObFNS/JERVUSQr0gmY
916hz1YAr8KfjbXMyosOZcG2WMCOaQALTlsbyLzb8j9GUY1aqrqqtgN2V+nXoveA96FOZH0I2Wbf
dKxvJh1ONjHoOMllhSTOpf81yul3VD8rfOJ/haroBKY52cD9/x/RiwcVfBfleWcrlX7znMA77+I7
7xC5vOdnY2ILkuYpXhe+evjin1wsQ3OUcOjuEArrJ9bFh3+JfExWLHIWvyyNsT8TX4M9jRFB94hf
E6uDmUfGI/Wb7L5NpeGZ7RrSSjdhfFyTedIg2SG1ma0mSjEeuRcfSJKv7Nqx0hfUrtEuec2GS67G
qlTgR/mOptyPM/t0O05Y2REKXQ1Ds58Qurafsm8d1OHfBP5/yg+oItYH+t1X5DSvng/9dyBZGHWR
yXrBjWwiVKwBwtVj1o1s6VuWTlMYEoXcHHCSoJpCQq6rxH5Gzp6xr/XegVLfdfMzXTigJtmnRjqv
5the6pFf/+TVcF6qz3Tcepml5SJHfTsh7XBWK0WaCJcNE9WJxNNEU4iMA57iT5ZFXrDPi2oeGiFK
Nt+NMt0ExeH7e7qKQuyOr3baNq1ONuWHdrbo/XJGapHU+yF7clqJ0gAgFBJ4/8SEifKn7/TzPdk4
VN4SjkISSs0t6iMNOEozQPB0/wCnfSbDnjw9hYTUU5RiApVoR64vdm3emR/B5NbbLGtFHWXcjB36
3CFvFo2jjIAIRF2aPmgV/lcjX9l20EBNVYnwRHzX94loUo1zUwTMOkrraB2FEUNTOrwoDas7+NbB
+bc8Y5+2GKJeL7BZalSBAppkmDpYzv7RpvyH40+ojbG0RvXZA4eZEJpUPNU8Ewm6Q02Zt5otcKM4
/m3Qo8nDneFpJwKLebL5gCyj9ySH+35g13LLT9EDXf6i4dvTje1YqF6NsvCUGwqSTocQYTqmzzVc
vKdBXc5Dc//odQKI9lwhKdrpnxrdKFnjHia5OC+Y7N350GYIXLEZyrvbNM/uenzZMVgzUbUdVSY7
f5wPoElpZXfTy5hi7U427pKwTW14uxmUQN8Elvz6tjmc9oUztuU7ZiHSibW7LsTurur174xoUp7A
0mMGNuHS6N4OQS1+8HzdVf+Le2ObTGS0o9do38EePyCv7Dpcm/quv+jjmuxcrmzoHSXPUVq0/npd
9kSR8fHOcfxuGiu6xIbzt/I5Ot1wOZWfjEUa2UKao2xK9RyKvhreki8l1yr6XzXh/U4rLZeeJpRg
0ZyfjvpIjCTy4jOAUEFb0m4kOjySDn0f5oFKrQ0+5NYOlL7Mag2gr4pm4VusOAN0ywBp75cLjvqg
XyFbiX7LYDomMbnvlKCgegsJOSoGrX1gtyvAu/aJzBHHROe7/VI3sBJ46Xs4SCrAG3sJ//Ysv0EP
9QTSkoIj5mo+eKd8QTfd0Futax5LTw63BT347fTu9Ax47FrmSPnYy4wlvH90qwawfYBXEEhffd72
J/wDLTKpxlvx2iY4XytAK/tggzCKRgbS6Pc4jOwQ+NLLR1QdOewetMLkMfRxnR1+IDiVgebO+/FF
J17a8w2+rb7+eEwG5JHntl8rwlQ5GRGSEvkf/PyqGksGRoGZ8KZZsUTwcfElu+r48MC0cOFFBha8
eTUGmNHBQnVJzmSb5KKK/6dzSf3bk2ny5sspTgu74pJGl2n9FsCPxzBNM19OSZq68TIUp8/CODZR
9LwF/KCLM7bhZVB0+OXGkBYo4J5wZrmHVTE5y/Eivd1uXwrt2sKYDRqVPY5Bf6pIUSUFIq/jCVW6
KX9eSQwRhGdrHwh4gFlDadGU/r50muAkIVjWfhru1pi7H+mjZ8DcBdQJy9Q8DmaNXNluHwrVwPtd
NrZ2FQ82M6Ub8jpFBr0zfen1p4IM0LpPrvCoPDDciwx9/I22JL2n0odvYw6Mw4GA4lzFu4Jyif5N
MagvQWl1g7fW5OcBG/OGHwMr62YjkQv5RTsfBtUhkX9Io+fBL/7aTKtcQkfOsgUXyNFBiF1LTkq+
DhvxkqJUnKFROuMJcZ/K7fstDgV24QSj90sOr6fUbhhG7oIpoPHeUHlTcl4rGHWKYgdmbYsSvtBn
XlWiBgzKHueufeKB0kvDjfqteEu9vNyqzy09KIgd8q4rgR2xp3CXnm7QdILGmzRNS40NLcKmUr8K
DZdxYzwpixJQTbm1YoTMpetdiESbutuotPNEQ+p0HBKNgUCWSgb8BF70Jtq8DfJHmMYnK+2QYc/3
oot8edPfJsjhRewZ3aNZBOckxZ5S4Xz9VqvxEQJuuqeq/pzDvIZ/Do2qmSrv8LFR27LyEWk6FfN+
dO830K8eG+Q0gdWRxx3wo0jQwzlQJFVYL9WMepm/c686f0CV4qlM47gjCQE5PZyLl6nxH/PWO0z/
M/1fPyTQJhXIWaD0e8YkP2pGlfe2iH0cyRxJRKuFe6NLtOaahJ2WaGW00zqBHrYeIqPtOE6XcXW7
z7SqvKJ+Lwd3l4rD8e3V87FGvLf15eKJL1G75wl1eupWnJGhC23Z27rtY80hAR0P1EI3X2IIhyqd
I3hBqQsu6SyyhSYzuKVGl3tvXLcmSsf7lKiac6iLI1GKx3i/VPX4Wk1zl95TdLG/z4HKW3tpIMgE
vMcP2mmtHf9mnu25zrc4l4u72gN1PWHnp99BJDPRIKjkn4t2TkJOW0BbZTPjzP5s8M9317bYhbnp
eYD4vd73RRu/YQF6sPCHxFec7wQG7rQniEKqd5Lfne/AUmnzyqFZnEHZfvSepaN9Llx9hOKw/tY3
Wc0tak38DQcYj1xy537dbSv3AptFCDZVw9xciFW+sMtN8op+Ajv5YYHp8KRFOV/RkV44H7zFN4Ig
EaBjxAvMPX9nswkCG+Vnyj1MTn6QrerlkFNpLMTpybltBowaqZWIwDQpNtkyz8Ucat1VbJucLt1U
wpRCdOkZfqsw4rynoYNqLPQYStFmr6BQ9+KmPrsK0wKtAeQhH5EvrbGeFrt5ba5LnBF8pFh1ecK0
X056Bkbv+OybdQ4d1etvJPna8r64MZ8Ru7UcGyugfklvSu4Tiw+vkrXf/WTA1XEhT0SJhFC0EdId
F0H8ooc0SegOEt5M/Zi+LssMh3B8HmbkHbv7uk6vC8GxzF/+wlYHJsGIj3md0x4Oc6nynzL2+bWk
rxI0ch8QabEprf32tbZsiZWSEs2hhDcEQzV2lWcTV6FQk0DO4NRTRJiiLJkdMj5m7QZt1BF/Lile
xCiJjpmzPcgarraovl4l3KHJzOCb4htEug8RMRCe0IkXHlxTloxMQzpHH80jfbPMcfTW9Do3EKlv
RegN4y+x4kmCPo6qQ7bjNrGhP/dZaetweMgqj1U7iJIJgSCzEAHRAf+w6Md77i8OXtba5wM6F2ex
N9gJqc6EMSf9ESqJt5q3jjtCpUL6EmhC9NEM5bypiefMQEt8d38H+Oz2HEZDWTtLmnFj/PtlvvlZ
pOOxMelhr7lhEhIPxQ8aBD5sdFVy8MetkvoCHVldtrkB4bBjLwZ91kF7mqk4L59ePynIfMUrUrMO
maKFoh8iVLjNhA2B6gdhAwJt8lp/zOAeUb3D22Q4pMpSOFcZQI2+GswT6DA6ZJjDwZ/rPoIv2Zvn
Y/59wtMkfSpKSKR40Ym8QjBFp6+eochqYTtXphg/qzwFOxgkms/X2LuTUmrCiJvO+hW4ennUGAOW
VhO1/Dy+cVdTiY3QLSl3jxfUFbFfsGWZsKIK4b+T8jeQ9u4/2lvP3Pra0d7z9NARq08O7uGVIId9
WNAQND2fNy2+7SmsvpiEbScGeMC1p2DTMaafVce/NUhXi9uDuy+AmOWiL2XzRIcwycdHRfnk/gCf
jNPibi/GyUME3Y28lI4OSeyx0dl+xqZB/sz5DnxeW6Uq5dknRm3We5WgMQJIihD7qh1I4Xmbr/Wu
qZf4EkJ8bOCdsG/T/CsXJmO4WqwmgNCfZzYMKUNFArgpEy9DpQrKtdNxHTrmLfH3JqwXJdjO0CF9
ff+SeHemuMdldSKfksD1Tw3VYgEu8klNGtRNIXy1ltMEnzo69MGmEGWpwlA4yANVsB782vMIoH2e
QORQ0kxT7dypiqLQGHUP2fqOuGq51IwgAjbjdFF4Ld2R/2nTd1h5PbtXtQglzlEE4eyeW2prKTGX
onKYeDhdhKSD7hM5972fH/YKVRlZ0iBjjg/o2ADGb4soAVgvAuWKFEXUFoCl5adBsaOhVQAlDeRO
cHsoPXYrr1u1Sp/a9z9ityCCazBvJ43LemZFmaIvyqgBAqNIsaJ3suZ553ZhLOURqOcO7Cwd3dWx
PRslGKqWzfpB92n3wH2nIojAZlWqCDIGSgg/A7R6YXWrjiabwM5fOmGiS+na+xTw51J0+bEXNNMP
UyLBNZrV3prqIBzD1r1zlxZXJ6RAkMyT4Ar3KRoSfur5KLuP6Rf+xHKucxL9+xKiWxo97cMd1b/G
S2pKmrifoH4NLc6yiuIODEs0wK3w91uIzx3aXQPyN2gRrs3/ECrN/Fqqi4yxBBDOE6ow7ovCnwoK
wWSVsqpxCPA9WBDMJnysTqCBSZmBQbTTS/hmG6ZwGVYZuT1oOHXTWHqdi0f1GivZnLvzV5fcbsVs
H5rdmQ4sjOzFhFWE3iU/tJwIB3WdbMo7MHR/yz3amYPsoT89tyyfCT5cxw2oT6ZhKRuaUmYP44HK
dT+bJanFboBNzvFXA8MwhjrA38EyvHHH5x4wJR8nJJ1keQJPE9nyYIMWI4vdUnW2CXzCXGiCU2Ku
6zls8img64KvBMSVfGaTdSpn8F4TEJEgiF2qk4dB549Dhp+btZf/+MXuF7BhWwC4lTQDlwg14r4h
pD4Uoy/4gkKgNALe0W9lyr9yS09+yQjLln8jmTf1sCXdeSgxYKd0XquKVLxeC12mPBcbegqr/Tsw
34/kSwSoodMtzedYlGq85hnuy3DIWqpdZ64ExJVadUZOiR1tXHfd5IwEDXCMbWjW3wwB61CqqezZ
VVHYYY/tYqiKabb8aahm8juQGWQUYM1w3SgJxhnZVbpXVcR2PkFVVK1Ct8LidhCt85ZBbk3Y2pa/
LDp7+bt1ML/UTpFt0tlZZpH/8Ba7ha3FY4/nGBMhEmNhIs4xUCanKaWXl7CslNl8axgfnUaXrEg3
sNdrkwvglSRneCYS4AbdCz43MjriDOJznh2YauE9XgJq5yAYsEGUwcmOWVk+l+HLhwz8sZE2A69B
pTwBsD9M3c4iujlKRsrOT0VEMiX++bbUwy6CFPu3dpPGaCM4b64jql+FcDFSuW8ITjsdymxZbXfd
HEUQ1RRREJ7SK497+p/PGtKkqW+YKpR7fdsgf0yqvEAqJ0byCdNz1b76RlAYwjdzNVtjfvwoBUr0
zsv6R/bkweZNZZTRjpevuQYDvKYzJsKQXO1UpopDAEOLpgk/ayu10GNpPx4i3bmo77n71rwQNPB/
5R9InlAgxwdnX/VkP62uDa4ipvz4szX1b4K7YESHHdL+3orDi0IUHP6ia/2qwh2sR2asyuWAqlR+
NR3GnBhPff3sxUECJgXfl3gq+FCtJls1FsrvWm5HUNc41vQoyxQPuQKohuR2h4kddBDFsZTbLtTJ
V9rwyvn/w7AVa4z38W76Rkbt5HYmBIcCMFaWhpkAehmTn7lHsspW+n+zT8dIZ+/vfzO8mue684EH
JH6srgJRQ6YtXHSeU6VvbnJphYK4H4d5qouQGtGPtalOdehK2YMXkLBzCsFb/wKMPfCUHFi71zpW
m5tlxdHc5g8Mk2ORJetRj+rKlwMyfiax11Mbprd4rZE5gUN7KdVYH6Xdcvui3p+26Kvf3ihsCJJG
u0fHsNtD/MQ1pvUxo3NWRVLKQ1yCiDxBM87rdigTIZv4+LhNE4NQlMdzGCf6uKo5vhPSIxrpLE2q
r1nXWMIG80AvZVYoa7TgQkYt8LO7kh+rjZymZZJVM4YEvc9JL4Vtz2QgSCpD5KbRYxorgSihlRNL
TyJApnUpwurmuxuLELKOva3P2qTFVEfAmrLwPBC2hS9gxgVErOWFqvV9B1yizq8l1y12fzxHewAO
UMGxhR03Xj864e3li8reLLS5+Aa6qb2oT3i/p4+ltJ5vubIa37LLCq91Ws8azKfUA+Wy52I4R9yq
QTyrKIdic5d20SRvG3eQ/RGumfvr6VAl6MjJZHzA3E2nmkm12ldBJ+A5bbGevXCCznCgP7FfGQ1x
lStazaVWaTUOK+ACP44lSI5ZmwHwKXPSZF4RpXly1/Md9406xVbgvTpmzwOwyohY48S2c534j74v
NKTMmJGeF/V46+fR4CoFgOseONYETs6fL9xUXoCXvrIHyFcQw4W2KFs/aeWmZrhJqGautNU/AnN7
MoiKkeeMth8p/UyCKo58xw6a3fVglbG8OZwn/i2VW+hUVN8rvCwmy7MqEGslyoBmbKrpfFpRoS1m
os55B4QBg0QGGoRizP/4j6v31lDF6zKrFBJvZBMBh98o88wBfObz62O4bQsHZyoEo0vatM31yIAn
HQigrIU1vEAEP14CoqB9FK4PiyRi127KnBB1o9fcsm5s2XYrJWA/US8VuYgKRHUoeibrqAfxLYZH
GBMbCqSgdnVJFLmwzWY6DzkRP7I6pMbeLQ/GjqU8/gL1NGaidHopq4VBAqI33kDhb5+XUckf+Urm
4+i1Y1NiwYjf/ktm+aQP1IEKwLfEQ3nH3LlLuWaOf6BihzuW76DCqc3YvxvOM3nHjyGH4NYYEble
A7vMZ9VmrqI5/nE8LiZ20aFcII3dJQzqQjr13Ja1HRKebC0Ge5PNrMHH4qm2N+ep6JxpS8EdH41j
E37w7nVJWjwKeFBWfl9PWpsui6PVVT+s9pRh0F4900MKxILSNFwtggWHor+jPRNAlX9kiUHexrOk
RusDleJd8Mv/VY/ihR+ua7SoXuGlwHU7XuZtOvFA2STURWfDK54fhAXFiTnFHlMAJ5bk1iDyyceI
7Y7oQwFWp7nKDnIzfMxvaqzwHAW58tZd3QZThXMMbfX1DMxMo88ezOZsGDXKytVM3BQXllJMRhkl
7FyEDtaI0PGCeZeK41WDtcE8IDQP/Th9cYJhBJnLqQUCQfyJ0DOhDS8j3bf5dEMtd1odM9y+Y9vY
EqU7wKUERg3B4jVGbYPGDZJ9pNodjbwWrs5l6FbhP88MAeN88OcD82HtYEbVl/Q/WmbESAxBJ0yv
R95ELZQBpHoYUnnIe9l876Ko0UdRYwEvo6ck+FKuReSzZIPmOchk/Y5zpNB86jZyJR/FKOWjeBW+
B5M8aAdsiVcSgQ9FhIlQ61KmDQ6brIP8Z/q33VtpXVSgEVUCtGc0Abvx8nvPUvNEs92Opp81JUQD
CdraWoc/OuPPZY9fN9ld9NRk+kvvrmOiWQSjzjK9tvXcOCSQjzK+M2rpe+sGDuNo4VWzmHsVbbpR
Fy9LJJGUTvljXwhybTmocM3UF230S7a0ndCXtskhFCS2eQEHd7sbOX6VBQ4xZs+SQ23AKm2CgkNS
scaaGeA8o91xVA+Ym8CjNsGwH4r5DDRRDdu1PHSsLcFkIwPczICVpOG875bGX61vZgU5QbfBauq3
fa/xLhYULFnfES9/8/Ey/8uilbgMc9EUsNwxlnPF78OIg1cChRRofB5cN0CN3wfBw56bxouhuKUb
QxDSySI4v8WD+j+F8zLDUpIvxuwRSyGi2KMTUZWFiJSde/DEdmR96ix9epscrcqLhCJvrvRZNaJo
wdTRsG4B24uErHS+QwsxTZXwGuM2+efo7F+m+nEZbEwvT4gS/kBxv/8jG9+SmVsm+H4KgRCwYJ9i
jTEVNC08Avril/rRbS51uB6e4VPbRe7dTafe38fXeBo6ATXOqlg8zCGWFb+dXKi0zrpd9FMP1IT5
u1EgMpaUDGw9FhFOnh1fNixWiH/YYME1hieubBH7i70lVPc2uNX5KOtHGZe++nEocZ7DrNuyOnc4
5J0QVD9BXjDJnn4g/8PYu0ed64dP8iZuuZaRK+L0/b//smVWN1zg6wqPDs1FLp7Trn255jjDMyx/
uXbiC0qXjOixOqRz/FPEStQzJPHoSoYvFrErCGkDKjmZOHy2Bk6EpWJvJYY61xmUr/QW1ugnn3JV
7+DpQ1xdQkSShAsGIBH58JzMXZMg8WLjn+uK2Vkz96GHIKjHPsFywqlTax0VUIdqQnAM7lEQzJqd
K+W3wmpSC95PSv68274y45BZ4y5hE3Y1xtw0UMsRKETyZ2tYTOFfbkH0vSlE4EITzrt/vBMP1JRN
HOwhZeHZ9wqOfDUAB7uLBAiXLtd/aQdAkipE9qFRdQW/7XOsp8LObkXg7J78WZihbdoak04eoXZ2
TZFKlb4CDZJKCF7oRFBFR6RekyygxyUet1tMxiOFTsQ9WiHaWugCAhY4HdENdrph0I288xWM7JEc
9+svFurkuyfOFqrOTXZTgbieKgSdQA2nmdslvltMsebYfuWFvY02hdmwfop1COf9+qJkpteX0zOe
yJLpOTADRY+i0QQvJ1X9a0uV9EJmhq+hMLkehZjj9nhPn7sIyXpET1sqF1waigbN6PO3vDTaowRa
xf5BgXwjVsg2kJ1TErqNbPXAoD24N2nL/UP6BBLUcxDizJXvHOjAdd9Vva/O3BGvBLjqFBTK4iDm
7ZKfAQQnLTi5XO34qX5a3c5c6GmgdPMRGFvfIfrDi4zmw9ebDvQHbdRysfDgL1K/F1B0I2vKBZD4
zo6OTQPF/INJig9Z4rpCrWf10aOV+rJlXzjh1zJyBH6bLMtFsxJ4ZuR3a8kH2/LkbGRT9PxeJZLL
HZJueDsCRrMJa+5STvJBFQUxuu8yvFbqTaj7y0qOLe4dOuN3WdT2o0GZ+qFnICxAQPQJmfFUTtTt
9pPNfdLCr3DAIu6utc+u+hs5OVGFObfiPSLYnSIT6redD/pNukFEEJsqwuF7LDrYH50gJEcEMXrA
EbqxwjKmXL063jYkMSRrYmGTTDh1Rooh82GivnR8aVhfmIIxf/qkDz1E2l684yPUWmdrp3+SFjct
lZsIBD38XZiUmimd52jcH/4I3A2sJpKQlaQwYRj2JJZNq9VIBRG9P2nvXWeJx/JW8g/s8tvYVWQb
MJ4HLYlHDSNwKOWRbIZxQAeNegsbdd25+eVuul9n+IT+LTG5VJFbEw7s5UtnSr+y43EMQME3cHW4
fq28+HJcV8En2Q9R763+ZpVan8EmQjIbPlqcUuzVGMjPQCd8yjDr8PrsL9TP+8nB2nTZdP8W1YJw
4UdsxY1l73CG6XyRFAiGpdF0P1X2mh1hhoNtR+P9l0GZG0EjhrTBZsdyervgxOSrRiAZB67svmrB
Xtf3j04pFV7wrdKPIcDMuBcK2b/A0XH1fr06hgFE1FiXxVFlmZ7FbMAzBIrXrpqBmi4h+bZkCdr5
hi+AjH1xfREIMtzcKGOKfp83fVVj/H62U6OgsA0mrisPSdhVjS6uZwJStXTGv/BPdsTxf67Q/QFa
st/I/RQrwp0O5tO/3WRsQ7yctLJIpfqihcA+TbISlMSq7NmTfUzJbJqfe6exRSM/fhY6nwuaNQdd
MY4X7H3tztgT8jybT8/CoS5jRNz9jOfSSFEWuuyoUhLjar/DUoJfiPRL+sg/dcIHG7K/+xFXLyp3
xtzGu9t/KAqEuUe9jG5vciD0v5ZK4qI5sZEohYCQbVtEGxF5WG/FKM4vOmLJLWjOOsfSXOfjcaH9
KCgulBoY0PTdOdtLYvifhMsLkddpg0Fw3lek+0ydjE/5UDs74IVFLw7RPGWotua/xuWlwe/kIZ0I
D4iTpw04IT33usHzQCdoo5A2fUGVxhv5h2PAk1AC4zYn+btWY/IrhhfKzM06arPNHFj9dHE5iG8h
910gAUMQggR5aLHIeACdRvsUJ7185DNUD1hPVBAbGG2oH12LnyoTm+Ca2po5onin95nk4IERVNSo
wVjLH2nbkxuCruarQJ/YSmFnulB1Mn+OaC1vzBrfa8QzOv+ABWFv56DKa9j/sPKVihtAYNFtzZXt
bUhQJCK4phEHowPlvbQw5X5Glr9KZWNEmsiSY3Fn3atz3ZgixtCRZ9HZDtfB0a/8G2z0+AHDyplw
i24zdRVXyyysYa1GO58Cjw9RYluroN+5n6SxmEeblh0qYCeVu+SZbZR81Z3ReO48kf+E5+ewynhF
InBKFE8aZ1AWLgntFsvJGOoM1QEZ/ciDtJ+ZcJjdpF9tVSPM5SZGEPdUsxjkD1Jl7recs4jzb3+C
OIw8AP05TCgfzrPllv4F/V4awmLfZRTX2aMO/JF6GPz/zT3byX+qxVgbMf5PBqJxDmlKfyARo9ms
N/xp90eJwdxKqcKTnPj3evoDf9AGuOCmvPoQulR6AX2UqgxG9Uwr83UUOiLFNtA2fbX2ZC/gzw8i
P/RM8TuLQfwwRVuWEc+sEjV7PTAu9l7pkKm8NhewULb7E2AccnO5EcITN6m7fwvUUkmfvl+lykO5
ljzmMwfpbD85H20C1KiARXnx3bL3fD1q5vuB79I+l8Uw7em+eCQDzQrjdxCURQpZvFYTAcCOl35u
5DXVnVEk2hgJxlZM6lFXCWcLJunR32ZfT09oq43vmOdqlzMCsVr63deHk87uFJZsTN7a4K4SNxFw
PWUImALDeVi2nh2p4gGOPhGpxapWfkvIFSqhyeQf4ZxVyetE8ThiJidjPahK+CQsT3HHxqHgyDjs
QePQpt1Y+xvQjDO+0AFWz7aFMm/VoTsxAJH7fZnSLj+5siVOgkMejC8ujnkuIsjUOp1BmH2yPfsf
j+ZGBG7t3yrwA6bIbayFPzmDcdwmjEAXVMeN134MgvnK66eVDAV70TEOpP51yVvRTvyx6d4M6z/J
svFycjicXdtckD2YsHgIFVoqz0KKfPIrlantrNU1nW5nQUku4a3J6Z2GRBAQCuaIylN+jeEW8eSy
YCxkIxiUqWOX50yVlnfhuNaqzzzl2GyewN3ZnmDvdyNzA5YwbbPYk1lIQ288BrMKIr9CmNFnVF4+
yug/svGVX6hVbAnXoizVKTZSLuFXbk3s0bnAVm9vN3AEeSnsSJwPSq/dUufq11xcLIfyjdImYka/
rNXv38ZNgE45ZP5nm/sWta9kD8xQAgQmyf7nHb/dGCLHX7dENKRkNy9gfwS1KPWOYBTJizneNvmB
q23FRTuEF/TkW4JshRUIG3zmUZYWaCQ7i1uidAYhb1q4iFz203MvnGRGPKhKcsF79ynfw4XobcTV
dnc6uOogmLFYU7H7ay03DCScyK2e37SXV0P2/9qHIcmYGenPdTQkDoAdRmkWHetFsv8vD+YDwh05
SUBxI6SZaGpGlNwONtzE7cL1RsOgBeLML5E8Z09znMlRxFasUWk6scgECxXnDW+wla9RiStx1pi1
zT773QnzOGwVmav+pl8LTkc6M7SVcjQTQjt0Z514WpJ37ru9/lE7m9xs0Xw2kgz2NlaJFsxvjyJv
bfOm4NQSNskUFoNhn7c8JT3wpHHhl2AFJrtdrj1It0ht1+9mvE0l8N9yp1zKfSjVTpCfjte4uXVy
ruKX1r9daAA1m+4RnEqxmlym1sVppz1OPH8ykeubkTsFRsI5LeaVWbDNg161Ri20rIx9jxuy23Ng
glRYbHR4UVUrVRQA+Dta9XtNGjic3g6SHC6k40/uNilMjA9ljF/0Eta0FGW2+m1peDGXylEMB+3t
PvbUrfl9y92UO0fqcDh3A+xLVcu1h0EOA45lpIe5BjquAOXnFKbOJnInL4uIGbrD/z9F1JmIqHIb
TWs0HmDxEysCnjbG4V/8SPfbqy0vkUgiCJsNu//p7AHO1K5Hl3v2zgKcp5ojMKdDcyiaQw+cf5lV
CfLHst6AhicoRUx0wWgadEmVVevqIa58r5tasuVbwyqXvePvEcd/xq4/VY13iNYbCQKDw1QNOsMD
jAkpMb0E7Z3q5oMnYp4tZr8QOVXU8DXzOBshmsyhFKAbmPzNwMThwUmDiVHjOHis7HUXhD1dbsDD
Zmr9Gn95iYLNmJry/UYjRq/0P+c0o9Op8J3vPZLQyay8t4Hn879I9nfJnt8KwiiahZp/Cv/s98F7
goS+q+vaLz+4Vg19W3hPw8KS630tPiowDi81LUqlk1WMtgTyPMVlae7SIKdZo56iwDxbrjHFlKKT
WoYOahcYJ4qXvAt3uZoSJbW5mJIEQ71A+d2ayILSZImK65Msy9s8J0mkIjjkCBp05ZUBPLK1yiEf
U8jkCtgTJ5IwS+DYgJ3mhAptW2e4fcqKqoXG0FN/XugVsfrTz0jxLryj3uMu7qXcrYD9dZ9UWnUe
Bf+cqqU3XbabCayheuHhShzxwLs9yEI5SNJbrcfJk9/UTVKN2mnhUSmfnXCLEDvVQ7nT1dlf14PP
f2NAh3Zz0vEi/jc0m/fORvc0U7MOuivZRF8aRm+UN3K+2OlRQogsNDUsqBN4x1Ee5s9ioHGZqUGv
oCNeq5VlBP0CHpUpQ0hyCmpuGEynC5uJamgiEnL62x06z/AVWO+tgH1Wy32Ckmf+c2Jd46TqeoaU
9Xynjkrh3z9pnpSLpsROzDXVWsA3ZAu0lUL0nrEYnk+llLvUbN3+kVDsDH32TROimy+l1/qIqgvX
nnvjYC5qabVlyYwvQ74ywa/FeZ+i5XtwNCD9ws8ffV+MHgv6b+iTUKACt10/aoQfWktjNTQ44Wvn
yX5QbSNMMzZJ1HxW95L9ZPxvRfXjBGmnAD1DGjQ5OBM+Jj2L7XL37nzF77AZTj5M2D7jTs/Uqr8g
J0dd7N+b3Nzy8WCjRZnrpQ+ebZnFZ8vNZzRGOTTH74L4lypdJ2uBazxHtZokUKpp/VeAV/3rBKTf
5aHwOok1XH+ksDM6LuHaFQyELthffw1Y5ICcqxcqs8RGPNT+e4wkPvUKCVslY9dQhu/IuTl65gDa
JPmtJYVNl/5/HmUCV0PMvYa1DA2yfbP3IxC3bBDaXnzRdHiA0HZ8AY9cekI2ysvNWBNnWX7cVApD
LnaZcMrnzxAgDkGlWpI05AoCtLUC9E8F2eUMjCxHZ5OO0jAuilqR4YgkoHQlGA6OlLYk4Lq00GeQ
yWRjuROSdxZ5eABG/6RUtMKdEUEtprhklaPH6X+alS96oqBs1B0wgr5uvU95vJ4SUGaetZO3UEMD
/8b46UwJ+tEYmHb0p4WiQYbokuSP13Nx+YTDWeEK3TjI9pC4L3bmuUCRC6hkra2ZLgcwPZoXPqHz
yH+gvRRYxn+boAR/QxLyHOPWTGyUXX1uS5jQZn1CmeEPA/ZphufBUBF9YFZWSkBbN3H+mJPJBs4W
bsYZ0cy0hBUQhhDMurh5XTzFYfIHHZNzzfsJ5i/imS949tusJslsfMDgzIlLv7l9D5gkvwhepuDX
4PL13BujpWrVoPW07oPcd60tgKgw9W+FLmHuVXDoQKy/3PQOy4jHtPs35IeS7CwFRV4dHSc228Nt
gNN4WqLjboeeMYCWoDwkvP9BWUhc0qp8MhFX7Z7iMGQBd+O7/i0m41XT9HFasEZYKm4Di4g7PKer
RWZBPURw8NB2xDds0ExDr6EKIkx6XN3b7JlepNVRLdlsVsbJ0dSKNNorwC3eHwsO2zavzRAy5qnO
QmS7QC6ZvXEJcrwgtWZ2DA3Ho4Q5khYzm0slhna/hMH0YkeBfF9JCoGp3XIGXfeZ+VO5D96q2UrU
QZihS+XL9f7ngHHFT3TfahhWKe6bLV/OiZ1sHcTlg9kVAF0dNQ8rapQrTkoVOEz0vLt1bvCnjUEm
DpiefhfSn+Xwe86amHCAW7AZPr7XmQ3HteBDMRGjnHPTTBvXSDRE7Hl0f5/kRdxGQUrx/zk17hn+
E9S3f7BnF7BjmK6kB8KN1KVn8VxCpvDUXdGQpSNn4cFUbucEn71eNw3WigoGyGiCCCbNaIboQW+U
IWMQTbU7Rps/MKCHtBBJ4alqcU98koQO51JbULauHcg9wdOvR1JArrMzaCdTfkKq+DyfkdUmZ2k9
03vwPk1fzhdRMnOjt20K//6zTFXq7NfHNjTwlHAtPMhPQIm6vqz20ba2Bnoxc9I1LjzX9HspyZIl
9DtTdBAzvIcG/p/W0Oy9eMnTg2Wo19SqS1oCHU8d3F+OzYiXCL9VGSq+ISCTxFwfkScWYOWpwwfn
p1f8W4NKwRDavP0DmarktPI/o+9eqIHqretHttp/opODh9pww4/ROL0Pp+9386tAbDEhwMwhZbOg
Ge1WL6Fk/Vc6EdzSWpkQYvNalcmxfRf+SlOy7RZweK+zykXBW2k5otgM8KiP3wbnCmH3xGLMNzom
7AY1xZCoBnxco80Dhq2Pzo4O/HRKzz7lT2MwoMtW8WjV/cdzR3VXvyKkKL5eIpHFGIUldQhQwtoE
Y7l5Z10Qi51f/5iUu1EWe6zPha7BN/du5eIdgL3zPaEQ46ow0rR7q3fW2T66ILPQHfshG65nJQ7d
xOBSSDQ+Jiczhf7ksjoOWqMzdugOZSWmVow44Bv2nmXgRN2QdcfQNeCa4JHcq1kTp9yw9TWFW28B
BPCZIzeBf9dqQpur781NuU/14CN/9b6XCljYXMhUm6gFaV6CK03byztVaEbtGqOIu47gKgs5jPhw
n835bOwN/ZNtlmJ/0ZuHG/Fr4lIGeOaX3jwIPM8ofL73mxegNOE48gk/BflcTed6Uiek8f/HdART
XUKvHUTAExnticP+I2RAai8+4M/P0UYAlXAuC8ATj5zFHcouBZlvDUtMIrF8U3q4H3tediR9SUu9
9waVJdUFO922V1Np8ax8QoosTJZNgH6pSYwUPxsQKczfGHGmNuXKyBorgeSeCfJg2dcJkq+F3rUE
Rn+ijDtQcra/q3tAfpu7vJClRylIylS5UUmz2IGWVax/Ti3FDtXW48cgNA1lCHn5qqlLpoyD3/Yf
Q65rk4PYAGIRc+byCkl4FC+M8H71UJy9EVc9sqgpOq82XZmlVc2IY5UQjUFAYHeaATp8gX8A6OEI
cxp0oc5U9DkB7JYufMjidGSjUQnS+Jh1DlQDeNuGSG5OW2z6yqeK1GPEgDbrp/8CFQ1kbCaMtIj+
QjcdVw+BfatTpju/J1gOQCBk5l0hzaFiVsucwvp7A8YvegfZvRVwiA6WyHoxDyWoLmu7nzq2ReXJ
y/CFA1oNd9XQgY3ARxg1TyvojvKLhe4T2CcnEEuKw2mS3SPRibrAPj98/lIl/CaSthq4lH3+O54R
NQ4y+pkw8sBl5N389genjpOxWcpW6kCX8/eUlMq5FBYBdmZ8d2tZXRtxrkdJRGW0drOCnK1P/Vw1
li9F3S45B0OwGb8YwvWWpp6G43uix9IzBn11KEcvRGyQKenK1RrsuWJ9p+BNB/Hn3lDCbj5UWThA
EzJrWuGg3VXsNXehOFFdYNo9kWXA1tmeLmuP7NjA+gBeL3/YT4BXgnG2NkOFTqGdv7WErjo91WMW
TijNU0pgzZhbQGK/MJslj+XhEJEvLGcW7D58nRzlJs6GisJCcQMK7MnhQSsktsE6UUhmPfTIXnhX
rePt4h2GE4X0ZcJt/rmdjNyuk2Blaoun6zhqf2rk7hI4Pfcxogob6SdlL68OeyDA2ethWffwgN7v
zEROf8Gs8ZSnk3NiUtwGc+YpvEGSsAYd7PA4i03672t8TuMOQhUS3Y+jw78bsuagvFZOGTcm6QaN
rZP1mArNUp6QgyF1Hbxg8GrbwTKFcYdzDUTw203QEK8sbfSw92uZ4zKi7+oyWzq37t+Ul1GnrEni
RbUntPa9bxWOYjvu37Zlf293+Avkz9CJAV3aRnA9A3humE6oKP7t+cBi7S+PMOopytIvw9IBh+X5
7yFiSEq8YGo+nC5Bo5HLXd8i98zaWArOOwzbrj5CZKGI6SFbhW9pi1yFYEa+4ViMTayOXAd7ZJ/0
DUzQTncEEt9fhg2B1EC0BizWqEJMVN1Pl/8qA1KiLa8wiEnkDqfVWX0E+YeQlJWUWMeSgB59pc0D
IKzBdLRiXzBU2SomYH6fHyx3qHO0Q9wxPAT64Ws2VQQISMk05anuBek/rC6aTVxb0hsNazhk/yMN
deHUaJJRtdbqt+qkjgdPgNxfILacVyo5ZXruCBSUSLk+m+LKYN70Q71LSjPsD1JIrswJ82IJtbDM
+8bkepwO4XLHWz/HFengkGfJeamozMeyag1fwdz4zuBEHPMUiZmSTScc7ARI6elMWYVrHZ9nBfof
gCBc+Fzm4KFx8hQ6He0V0KactkFM1B4FX07s/kSbXkwf2hnX7U48nmzRCZFs8A3+G92BGaTxRRGu
F9AUDQODuSnXWS+NbRQ68kSyGwWyFL+l5OVHlwPiPIQQQH/rpi6Nwu2htbyoh+H29THIH4UubD8z
ul4T+ce/y0/iJcDbeLfNaJBaFrYGfxkbP2G648AXMZ0xAE/sVrMw6y61pmIQOVpw3Ct/Qb3cz+Cz
3tahflmrmMgAbW+O4h+ldpYEu1M8ndW9ncdBEHSC4BlMCcf+2B9F5QrOIfuHUa9/FEVROjGOr2aN
Vis+1eguvjYVYnPoxOZKNUaLu+qX+ujbO3nKQ4PO2NwddNykvtjY4CuEeZtS8MyOpItFRCydAhqg
VrjsFDIXYNfgNg+661ob3kcbXQ0GFPWVyuOVjgpf2W0j8a5r8jyHiUv7P9KblZHqKkaWK8uokShR
Mjn1tIM5JuBJL0JGluyOFis8d1vULPLfhjhD2kBDqFFOoPVdhsejDIxr6Kluwk2F+rDcBqvKlUlJ
YP2Q8arOKC+jXiwcu7oxrDOZq1LtOi1ekZjiVTLnYsr+Hv4pWqCusCptxu0Hdqfz7tMmsd+wL7V2
Pb3y3mr6cXtpF1ySL14JhUBeexNi6Pb+N9KXEZIBbyAyC+hY9DbG+CYvPSWfjiHl8FsL8JN6cick
gwUJ2MBmUTzLWq0VxWXOwZRC7Ig9yI3TlWmnuo71GZf7CcKawDh1ThK5/WpDOtugBbOjostr/IbD
aWZGCwPD/hZY9wIkdPZCYdH5F2bvYsL78GbWmpOHyfGoGvPA1MqMQ+DHEcvRunr6lNGaOBBGQV3E
3OInGk3grh2ZxdD15LO2cTomyWgct3piRvQ0vMi3tbEmsgRru0H3Pon2tGGBgOiz3J/MQPB6PCDd
jlnODWO9lSsE/2PZgweud907UBaFDhKpkTQIPKlnpDZq2drR0ntG+jT9LxAUCylTTu5jgXk3/kEU
o8YBMvZSYNM72hlGmBaeO1SS18HhWp3mrym4zIX+JZRytN7KzzfemYapTyVU6416cVqzQICex+2S
EhnsovhoQDs/OCRrJRDnqFTA/fwle0y30G5z/Nnu31bEqkbxWWdGxwDQfNu8hzqUemOY0egUh38C
/WPeEzG6BxTMJ66nVn63ystRW+b7oWfZN2JVRRcc2PUGn6kiJ7mstabMTfpScRYLUgK9Xb9a125Z
4rCxcvdExgB0Pig1w3Nu4da/qHW2ymQf0Fq/B7DqAao8w6dzU08FYA0NAdPruAid2XldOY7OZcVp
R1yGdazFZn5Hu9jq2qlc4txxkjjLsZiFsmrB3zm1XleYKlreKsgAcU5jXbQGRwLwvxIpv584kjvs
Fe9XEd1L2labHC5tLTCicHIZnic5XRH82u/ilriDhDWgv8z4njcNJSv4URMZ6FHrdvq6HQh7YLGr
9jqqNO5tY53iO4fXZWLUB/XSob0293Qbl3drD0r9p26RP9xDirFlcUxxsHWrUYl0Yl79a/K0R0Pu
oL2SKAKT8zJhxmBLeTpzdWKRB6XwNdRaHaXB7HmmKVgmpbZuYp2sf9h61n28Y0aKNROX/7YvGO1E
eLp/CXjQ6x145FAVxJQqFx7u6WHFTjvKUcIVMmjUnBjGQP+qBQPRkdW735t411F4w6geIKfg+XNH
aQvsCm3i6pUyu4dLoDHTbOGPOa2V29o0i90ptaeArgbcTczN7cgcbjoiX2UW+83UjMhXLvTJDkdD
QexSkYwRQVGZqnWUxC7yBdziDcQvSc9hQCEGthZKMAdsgRX8VYPPv8RwhDHgapkKMpeunDaJqD8P
zwWD6zcJD+pmyDW7Keo1L3IjQMeIvvFqJDNqrZb8UMSsVSfErudKyFasDyZ10Ob1iEETm1B6sEo7
26/NZmvyPc/ihrW3ArZvcbZIiX+lcUUNGy+qJaOoTwfjxBvmTotoDUBLPjR+3IAnRHFPEG9dLYnG
AeKUn3Dg8oio9k8mbt5exuXkri59wS9ncOITk7ISlahP0iWcsfOtYWcyxBWtNL7AxXyvryBPEob2
q8PAoVzt6+D4iANuNpiIP5sjFpqqIis/JKqmc144wgGFc5kDO1ZSrVIuIyLdJs4RKvnBp5GwtyRu
3Q8Y1VEND4pkM0ziFThdvRlfBRth1hwOKYDUguaUbxeJNGGGdzQhjW+54HZPDMqj1czk2QIvopB0
T/BonvpIeUIpvpipqhEISBT92hFNptHhN8bVCvIU8aAIBNb4STzlThdE3l0E8gDZiquqCadtuAao
7iEhb5BnTHK4L9aL/qZZNhgaRNkWpZgMeY8Poqp5fgubaMz7kXJToUT9BrnoTQMlGaFQ0c7/nobM
hLqg1k0V11fEK6ODGxfJSOFSZEvZ/WaMJxX3GmzhYOo21txxYUM/7gBythqwr5IY/L4iaWM3Wpf0
zwr0iFiJunq4Sz1R7235D0ELx/bCGp34VlXLpyt1EPMTMcHmVkzOKBCDXTf/bn7tIUesSU4l7gcy
46PJ+DK3xrmzR//20yYUlyvo3v9LDaU+tlKTVPPPHT5BjUChFwZ5xP75XJvX8VMK4qjES/VxOySz
KHr/6mbwgPS4bVwWi79pI+Yeq5QMY3dd7cluwMppkH0veC9z9tRNNFz8cWJ4CAUDJA/7Ikwl2EHv
/9reFBZ7tUJNGB4i15KCiaJjc080Yf9TghUdzRUNHf0tMDIwGtxgbJWb/DqBHxvEmFRuGFB2vlU6
bpSJSMZm+jHREkmHiesNeLlu+tbBbWGbN8NAwXza/W8ViAjq00OL0MyKbc+8QhTOGYAg4v4BRmOB
FdXFW/H845/Fd74lkiLSGT4ThVjjsDLRM+sLJ4fVkUS3Skxyhpt0MmvbSLI5M9YTJmWNiGmbhlni
T5dAWhFpZ607zJMKlkRMjBX2wE9cnyKMf5inRYOPsqlK3flhuTOkFm6nin+/n1R3Yi5YC/Z8DKOz
wd+/GQWx9iG4NTsT5yF6Nm/HwE+7YZqc/3hrJEm/eklxuV55OvU+PK8CEouu4Hx2EZLAS1usws/4
p0PGbehVPweweFi+qmhvcF1Ky+qow9P0/at2L7Oht7zG4Tr9RTEML7Il1vnxKKZdHWDLWSY9Btb3
m0mPzgm6QhTSq1+AGQFX3I3prIYGOe92jNaJmuidxWIYBB9/8GNRnrSnfer4tAnboiil2+yWIOIw
Nko9MCkkmmyZeTA6WVFzZwtKKClx9gUZH7aDEG3sqGN6bG35b01CCFrjsgOuYbwx/3oY3o28WaEx
5t9sLwxXK2KqjqHaiHvfEaaENrvSlbjgggP+pnbHYXsoRoPrRSRqngNw41R0XVGbwGtdofor76Z3
18xIEsXJa8Bq6SbPDskT4tM6sHBlFIB8CKi2a3ZlLsG6kH3H2dYx02Quw2B6EfocK6/nJ3pLE5dt
CJFzkyuf5Mu0jMJcEzeAdZDHLn2sltAnA3LJMhxS7l7dA21neCJYJy71YzuTRDtnyPdvIzjm/Cu0
tjvgg9nNeLLMQdsFYYmYm2fZ7C9PIGak83gccMlUhMVLWUgOiAwXIqqia25B5TX58Kwjo4QKy1My
TxgRTyMkq5YvTjTCCKCsh9t3rNlNDUiBYt8ZCjWLOF/vbX3pCflj24tZMStvk4QK16+clzuED8vN
LM8K/bNu/xja5yKgiiHr0O5xcHwqGypIJNWLUVtF8MIm6EHVDMj12CzPQ9GQWB0SA/QVvu/HXJhJ
rXvBPqX8gGi/Nsqv5wPY6acVcK19V63JcivVUemGaP5qqjqzr4s8OFKFZlNW4HSMnwfpduCRu2I4
I18W5TrXNI4aZyGKFeC8oVaA2YaWO4jrvXE897g//+AnpFL8L44O7Ch2kVqjLtmuJzPNSYPZNHr/
Iv62OZaTwEK2gSacslwOAH9RVPPC/Jal3b41py5yUN4vmofsBJZIDk8ka4GVCnc+ERKcwcXfZEp7
uSSz6rSKQCa9PtFmn6af7pHvH4VnS/iUv3+PdNNhvBez2Bagnq9b1Y2/yzFgQQk5WU6EIzT7Axib
j358lZntT4pNZhe7zfvubRLZNfjjGZgyd1F0tybQnkLByKp41Xh0vJxIThe4RynpZTXni7CqLB1X
naldhwJPXeBedOlCecYE+7mtyHU61+aNvG6fc+D+N8gSZXSgaYS4rS1hp/+kFR3LAqVa43WKFaH5
a9+cvpww9SHTTMe/4TwbM0TF5DCm5ADH9ltcpsR0tAQjgbZgD4Jh2x6rquKPCiQ7vebHOKWnhYiN
wlmyblG9NeDvqB0FcceCg3LsPnT2clneDzHKCDyGUx6m5vx1m5OsxLFMla9Nb+Wbxb2iXWj/mI6q
npf9H6lfkMlMVvwR8ChoJHYsHbjaJ3s1JnC5DXqC2CbvnaKu0qziwS3BqtKBImqJXUhJDdCFypHc
goGpJAiMwi+m00hej+VXRVhIkSNSJofcwW7eIAfKXw7XTWLabPD2WTkAouZX92LKpJ4IPfnnG+gc
gRxtpFznlTZihebw2WC7+eZZrzGNOnNn2CPw2/jKFzL5EKBTGUccCOhspI9QYGwONWnvcf2qcdaq
UeHV3C6bzHpOjqQM6naUrVDpAAdJ9R/GLtj9nWzhKaEy/3tomjKxEi4bs2FNlTeDNiZYDq+FWZL6
6Hfd6iUQrKtsvkSSUexiWdvLasFFlrqcKNW/GrO3OoL1HfD19T5X/3XKDVIQw3si0Bk3XMoyuTPl
P7IfjDZeg1H1jhlDVMNJaOdPLatPsXYyDEMLL8zRXBuOEdurgpw/lcamfLT/5adjUqioycagoR27
ZL5vPYh6K/ygKIK2yZdnGETKoBTCqJ0ukO/H7GNf8HN5vzdOi7KhIi5g/Wa/N/nrZTbbF4qkq75S
91HbVLTT1/UNkLfOOQ4u8AbkBycb5YHUDl0gftFWoHM5XWR8wwt2aTUphFHBJ2wSb7Mc+2UYpN90
eUzRxeJ77VHlylyQObzS3XYgAyRhS7p7sI16vOaTAfDE6G4KuWrbSVcu0yP4/bwwIOKtnS8P6ROd
DaL7EFnRBhOzjaKe7BYW95KIX0l3onav/EW1DpRHHaguriS8LBxfqXNYrw6M01mQ/iLjVAh3NgDg
7Ani/1Z+hluNjlfbOG7d1RGdGW26zxwVJWLS3HLEEdTw8TMwoy2MAOdYpkCHiiVGpZTSAfBDKm2N
czSA30994ESAaloEKXtngG7/W0HR3T3OSF/OUMCyzJOU6aaLZ04O2ReyHuN2nDmYNM2M0iu9H4cO
rDNgMBRgT/4b/yDoO3dbnz2iL9UKuj+rU743aae4NDRwGD9+3gf3ldG5vJ411n643EJtKJvEwkeE
cO/AmIglwVy1eFu+qqlxt1qukf2sjDFO7OvXDAdEdMmkcv9IS6NWHJBiaruA4wXvjpUHd8bMRh77
ijYlcABp7uRD8j4aJNGvu4pn9YPwtMBK5lz3fVGGxi4jV4wVhR24tagUQle+i/Foci/ITfdmIkwd
RGE3UA3IsKMOpD/r1LTbNwPuE1h7Rp+4m583hDS/FBV+SDyoiJanQxozfspW3lHCUEcpojZp4GCd
3YXlkqBCVjEhBGJoT7eBJcBKbzj6htfq3W7Mt9EsQBVQAJmhRppkqGkI6Fvu/nYkJCNZncXRKjeP
FtYEMSCSj5dPxNsVmsQqUJS3G0UQ8yIhuYINLnTsqhPHiZnmR29h3lQIGonDaKCFDqGN7GMU1Daa
Y7X0FqYuTLnpbgPUxs3QUBQKIJx+1+4yrqRV0gihdX9cKMOmy4gnUnaNIIcQHR3ILfUDXTvmdrrt
AulEdC7RXP8WhqAD2FL3i0KKiRrm0loCTwaiROqdIjDSu98eEislfezOxaL8NyXzDEIW00LYUOUS
KkvDFndHo2sFYsT4u7/eqwy0diQJeWlfhwBFRjJ2XpRokconVsf6ztN08BsVAByfrCtlPqnHMMf+
wimYR+bWtLxF1x+/0aAg3FlwINDgupagSgAnClGYHMMm2fyr4//8X3snOt72MIGkWmi+i0pjkEPF
xaU47QR90lFKzXs9ubIyrPIUqEO3cg60r+doWbWQGAt12sxAgHO9ksQ8aAUfMRC59TUXYXOyZb8/
TLvRDVx10V79NBDeX/nCP6w5gXD6Q8dMXf0mg2W2VDUhxPcykv0GRcnNwENJ+AR5ovGXKupTEjXk
vgiApBbdnmurzxlcqBdouWlPfW24jrkR2rN1N7suCBRqOwE7MFy7XVeLLAk6Nxo03RfIWD5vl2J8
dDbk9uDRlSBfK7F0go87klnXhBSFVlFx0Bwc17LLu3z+7CDDeyiD95ykEYE2hVVIX+yO5mfjbZ3G
gQWRga+ZUNGirExJy8TY9SOsQeMaa8J1+jUrEGuNWYzVm80Z/Sk4LDyYiD48j/ckuttu5Jax+92J
htTKxqGqohkm5Vqp6usKavLwhPF8YThybcLKtchcbSZaOugooRbCFHSnDGLNSKo4PMKwGMeN1bA5
x6NEBmodHYzgn038Ax9F1eUaf1NDMN4EEpBQP+GbnUVy6tzzttuEk7c63qGztGeaDyhhAjdIAUQy
Dmpe69isSR7/SjujwqtVNN1lqu41ndaKD7CwmJr8isU7kAJwHgGjCy5+rTDGOyjM40RcvQCGZqfx
HxZtqeGuq5OrlJh1UWw+b6v2RqaRUr2jFmB8hDcS9YInMdtFzMjfzRCq7jyecM+xmpxBLEuRRAxG
KeHNhjsF8EGquq1JkLfrpgaLT4BpQgkGnkhRwvfj1z3HwB/CgRFogGLsyLTYVyrxiFd1lUb+Rqyx
/XZDUCZSe0bB148Oc51BhvXFHUC/wWkEq6wysKISajgfuR629sMPuffsxOvKZg6jUGMrGceb0Xi1
nbb6mZFaO9FOpycuNABZuBY0dvENMivNzz1CIKpmX04dlTgSwHuIl10IH0hYad144lN/4dT7vcbD
gaXkH2u9X722859TWTBSK0XuEyWe2t0F8skcXSwwK/H/cqi2JRIhYAJaANfNMkZLQBeswgHTxL+e
nyiXwx+9WCu+VZusWDN/jcEs57if/O1UMeqkdQve7A7toG+uexpCiaXM939nXT0MkzNTIVOKXQ0+
NZTBHT2J2uOhCXOIQKEB5k2/JSLC30Y8jbrB75+tyi/CQFwbsMzwdbI1cSe2wzT85B4mi+4o30Mg
2QQmemBEwSUWwoHP0GopFwBf8A2TrACCobWN15foHpOFwMkGP0jVVEiBlWi/TQTKcVUBu9csLOAP
cBizdmncT5qM90FWqrGJssrRfiQKeslcXnTTREVX4TP4dS3R+WbrPzS7HlZjTxdiSH3FAzodJtRx
9qBZfC97+Ak9Lrhex0VD4fdDH/It20e1AefGNMbmrO58XT9QA0FcrABJrrgzKOZSizFS73ObrJlU
2EPhawW8sgbkdw6WZmyC7lWP0aJi2/PGRRIR0FDxnTRRZMBAJk7WGqNCuoxS2zMfSDVsBVNnQmXb
6f150opiy2eYPhZHQWxACiYggNkfgaeyF7c1HcMZo2+/Ep3T/sAOzhq1HSDyzndr/ksiXQkTRVfL
vwhJT0t/PZGNU0L5O8HaoAaHb+5AEpijZfE0ivt+DUTSLomjUyfhC/sN9gMT2Ki+hyvvOeIezLYU
MN34dKXGYczZ7EUXRrq8Oua7oGolg2tZT7JEJl/4GJDFYlxtxz/RYFjL/4KTfPWsQZA7LRrpPibE
gj8WijbjlWbzudBCVle8acdrzWoHy4g/tdjbc2LzfGQAPkqAVM3KJUESCo7QbVWERINoY8pIlPcK
LKcdsU9kHwFrbyLIYtBqINZqxnFc/O5S8bAknbFT+3idGM9pvACorqFWlLOWN6YD9jFMSkwqTLHA
PQlyVWLBPwmzWmCp7Z35fRn/AjIwBIPDeLTiMVm4g7V7eOffdbNm6IOV5W9/eBusQ+kcSYxaqoM/
hxwdrdADz64fqpP+FiWaYPHXSZ2acwCz9BltDIe1CTYilZSBTgWgVEiNhKtXNStlxfLn/xQYTuQL
Coqf/WqKZoeIjX5FRn2FT+6PJWm63mOdTiMvNpNXYXO0WF/MFqTZVLexbVpmjV6LLxK2Mi2jxoOY
7LvH1kfnQ/EuD9YEtBqvBZvvIgrobB4oUXnVqGsNoVtwaWWPF6LoGIIkfNDmW14KSjf4q1nbADjx
Yvexo/jBGgSMcB1tlZxbSANHPIrTCZ6k7clRT/6zPnaB3VJMW2BhOqrc0KKB7WeMQ16tmUd+drnH
ss5G8dC2wSUrZJ3ilVQcstW0UdPopTF7rJaeOEVd7YsQWxZWc34ACbj0pQlZk2xVfuVqrzqg/9gE
4/0LGjoDwDdZLSNi+nDp+ZHoxfHsVAeoI9QqRTNJ2nFSNiL3P1AMc3y6DUDT+zmE9KTsHbkW32Og
+UeNAItWTrC45xfSfH0WFcSbVcJD9oHyy1X9nKhio2HNjeZO8Y2G4yu5Ehib9lyhcIDefotIC5ZE
xWFDm9z8279mYsTCfDLne5/GyYKPhG3MR5Z95LZhGbVyEWc4P2Hw1rS0jmx9ArIoBw1cgxMjZhIP
9kgU9OmSJhmFL9m9TEAOg4ehtGCn4jr5iKw8DJbd2HUhNUVKhgkKU8LUhoArOxH2aeoge/FIUSIc
juV4CDInBhbr++41ZkrWrNEbZFFl0zOY6cl3Tr6XHakfDTiFcsWj0tCdJQUHfUMZAvF7cj6VkI7v
QHeD+X1CkY89xwxCaiaEeZ7BmHFcRStUNDFQ+5btnnMwnRP/Ba28y8kzN/ILmDMHqWUMv95K+tTZ
qNezjYSoh9AeaKJ4lmdSX8SX2EPOzc0FahVuubRbu2kmcnjwwjNfV8oYYImNb8zZjMQ09pRQkBTr
6EZzFqeM4z5FaYT6+K27jAh5neqFSrWLgL0ChSm3InYKKEUTxXMUOL5JC3Xq66PtXoFYMJS+js+9
+hf0CiBLKkafWWCZTXjJxN56OfhFfZ+KxT60hC8VYS8lF7Jfnr64eoBGgI1nD6dsAR4tVqryq96C
n2XKuu6eWFyKLiNbVhx7mqiIoRvoJoO4waAjN2uHOk2T25nuWpviI+y19gp/Zgv4k48gJA3D3cqJ
QFXjuzTsrhv9zWFBbzZeFw2PsfxQaxNWnovUywonJ88i5LoGfztzs6DiKwYSch9cw7kkHEJp0LaZ
C8qeaAeJTmBG+Suy7RyWlwEIPPkrdgR1+6tSrx84f6sbYIBlgHRVQFgTs3eV/oi7nb4vBcHqUuM1
QOt5trHTweP3whsBUB/n/UZ+ZdJaZ+bGdO/7SunXw+lNVQe0SXrowOt50lJTcApRRz2l4jixYEjq
BXBHZBB9NhAtuCvP5F2zLLKA7lqfTg0iZZc2wE06SHy5JQEcoPTSAxCyBSOUHD3cMmD3HfdkAczG
BjrYrmr3UH3lGRxIV3f1s8niSp7pRZIHgWz/7baw3OLelcavUXkrNhUKCoF4+zHr+1DBPZtH6dvR
ZJw4EZjfx87Mo7pyu+uvR9MEFQSYNS189FqIRI8SSxuhfT7qrPOUeuBgAS64iOFrCsPrzdHq6dNI
jfiWahWKnd7zqZA5rL5FfdIu485ASfODAhYSW77aHC0Ba0tw5EMX0poWGWBpFgckXIlVxOxaRu/R
VI6TaJvR/HaL1fOcp18ruUi8bO/9/Ri9EvtqXcmfpDj8tfskNpo9pVfrP91HWhHXNFbkqzwndFe9
P6LAnBLjDJ0/qN5W6mQOmQr5d/DRKeZSiyz9mgcuLTXcKHaA1oZHIz3MeEHb8FlUhMaIt2g2HLR+
FVQO4YtWpVWtOdIzfQFSmpq4iwOBa8JWQOnJNwSe2/8NuZv1WvPmx0hoC8CMPCYHaCKo+T5k1X1U
vUa6eIOtSbeIhBTdp+LMA4k0QXW0+YBXkUOnJTnFPTDdFqEf15TSKMjyi3fAkM1hMIKWk9xyW4y1
gPkRyHw5gXVBIQAjVpD6ZtZr8f2mmDPHn1sEgC0twu7eW63qHL6C+kshmCM8FBHcoquoD/QuFCBb
z1OwSf4Z4MSCAXOjTgbNxi1wTeNGoia0Tma9zknTwv+B1LR+jx0/7oms+2jAex8/0dG8GF6qj9TB
KjYNG54ZsIbmX9zEBErF0CDiOAc1106x8NW9za+s5mtz1Hvjcng6QUj47fqORcnGseqOlQ6uE3AL
8y8oc0XIiLilppzfmf7kdQo90RibTzAAL97YBp9dd1c12sADfm1qPDPz3NrS4NIqoseEo1t/3YVG
c4QGZC3lplFQhsO9/XY+8sYpmQA17IerAncb1m/lGIFC510DKSRAp/cpqmDLLpN90h9Ap5kUVd/u
/78VJHCGx+Bu2uHZDVezVM2CUCMkJInB25cczSOibb/CiLIuuywC438/s5h+N5leRpNQeKyrwicB
hQq4Ok+s/w9vG5s1CtX67JX1kF+k1iUMIw0JNDLPiDsOdKrIlQNMjGtIeT1OaY5Ku+2pAxsJbipr
pvaYZ276lWxSXSLqwHQkx3ZzJs4GTIlkDQPcN7L9C4UwjNICYAkXawxUiBZx1yeGbsIoKhcZyV2O
ZQGfRwXA1CsQIqD84wlXBBQqwNB++BdRulsF/SlUxz9Je6H7N3TezjltR9ixKvg220brWc37gcaw
cEUepPNaZ1b31TXSJ2gqdmQzb4MlMHDBDanv/79zOFC/h7YunOoN8RUdqt2qCGwWq3WBAKuSN4WP
Y0neFknBg4DgtYVzinZvQTc6f4CL+YYbY5PQK1BuRvyOn2u9xjRCU7dNJjHseW1jEmTdEhGIFKGB
BH9tRhCd013p6AbLvd6F2cxwfW9XCeu66W5rrMenRvPgfugtZ2R/pqzYkq6YANu7J8lo0NVF2S+n
7dfqswf7jPsn7RUgFYQUGBate+/Add5q5MPwQjm99hkgUo4oCjeNlLmzDiIvTNWuRzMkXYJ7yD9u
RLILEIQL4VIwH8k/aWcfLqSA2Z0XhBezLq+p/JfL5M6nptU7w8k3WTlXH+dumQhsr0TDHZfIvRRD
6v1gysjflRHogj8uw6XtjikbnQ09i1q27+yNDtQ5kM80DX8ZSQPqpfPiOSHTSdnIf7sUtN550jTU
kcJdKqf4GKGFzk9uGsm3xGe4j+c9qPgGcd1y4pQn08sgXRQFbMrFn0cB7tx8oESJDEUXXl5i2Aep
FjWIN79hoGp2Erfm9U/v80VwVhCTZoy+CL/0GrFDT1gSSswA2d0FS0Od+9Md3+7fd2xl4z+FqpGk
FKcdYvGfCM7d+Ht65Oub3614xTG+wpILUgmI6Xi2IiXyCyR/+41dxYN/XVtEaKZKfcONhZFWuNaq
hWKefwyiBj0x7hHt+P2Oh6QZlFFN7uAbI4qWUnIJTieDlb+KqTJ9k3gTOxZBnFYB4TqHecVtgeAD
bD7ptvP+GTjYXgtUEtkpSOJ5SybIizHu8G4vuiZ3Cx7U4gFAUBGV7ShIDza+xmLSKW8SboDMYkKd
9fgnvMPIz1RmMFv6e/W9amfZCo8pcY2NxlnG0ybGcSov8S5GXq6AwSm7+6jRaaCTdgcv86RJBH1d
NnOSBjHBviD31FGZxLapqfu8yk8RzeMhCt4BFbjFPO/zwBmODqUSOqkqWo4dPYyfMy8RtA/0bKXa
KpYwaUMfvl61I2wVkPe7gkP4bxNfuhn1cR4vkNf4pLNTxSVIgYri44HKBGeTxJcNtr3+EC+3RIgr
EKLG3ZVxYun4XgS9J9zXUiyiNb+Ab9bkgxD3IWDBlVuRc65KC6ylvqvRDX77yPpx3MzJw67q8PtN
M6tNpeG91NU//tARmjWRGZ08o5fFO7rpVKmRpX0c06eaJS9aSTmHkZBHm3cWQ1INE9ysdXTipBeC
kkyU1M8tC4CRx7ZO97sU3fxPmUJyLcubdRqlLUu8vsVRiKBKf3FEbeT+aXpGcCAiYdEcISOIXo31
+4Z5jd5r4M3nvEta0fdLXAkZjZqLY6J8dK+uq4rJwtTyj878F7PGgkNvzzruXJRseZXBl3HEoQOx
OI02zx9LhEq5AGKvw61P33qHV0X4J4O64cfddaICI46e2u9byMsPfYLq+VaQyFKnk2OJBFVi/gnc
iZpbPBnfRZXKwCqrQdFPXa11VtFWoQE7YwvHGuBiiGojMorO71IlgbLJ4ZR9op4Zsc3zeqdonTid
qmhm4X5n8lvHdmEAMhUvtDpHj9dW/NQbIvpVuDQOQPKt5oadDFzQ1ALBHHIuFwOEuPDJBvr3xKtC
VhCyJOhOUYD2wo4XpaBpQfc4yEVNFZYEJjHLyZjv3I/zvadQQ5gy0treJ4hPjNWVGJElSGVed51I
lYW7VyfJVurCHH4qY5yTcB7vH07KfDOxkTc0+RAaM0LHOZXm8BDDBdwJyJ2M3qLE9gm1rbZjABtg
doo61trfDVkEpsvYExrbzZM7YSbqG4IEZxX20as0VvgovJuqy+ChV7R/D5jdbPQ3UVV/6okWUf4a
71Cy5Vhrw6rrN/0xhE/dtFKgM5GQJhT/uKQ8BqStVMJ7xu7V0DDOSu346YuCZtH5hAhloJ17pI1f
dARPdq2auGixljZl2aPxRHDhg0J5mbL+Pv1zs52oIX3r1i5jb0ebTlGkFxuhmNtYme+M/yMJX1f2
0oh6m0zSX0Wkv5f97E9QRtO9DmGLZCcprrgg8xM3TRRtfIoCgTmjSj5kVrJUdI9wYn8z1r+uzsfR
NRiaJuzNAZXBmTkFqOhLzDwU/OE+WPMtChDPg1GABBvAbGwTiCRQl8m6XQDsA8Nn34VTLWifdAN2
G90iRn6JFDot2z/iBsY2+UA2WRUtzIT6tonjOIFHrLgGNrXpXZ1Bxnm6tMLKKtyP5yR5Ho4fqVUR
isRu6zZNMnsnWY8JtoQtmyGMjtbOyLZrICbkTYprC6p9fxDFW7CKlDR0SqCB1WOyynyA4OlH4Tcr
o/Gd7PYkLMPACUrbAlE7J+I7ma0Sk0jWIPOsndpDeH62a1cw7vk336unMPnVFN4S0ybwvYeGO6Xu
qGq/rGeuiax2Cn5QQgOesssIVwbb8qMqtWzRa2upArVmNyzoefGGtfZzCtJawxfwQd2X61U8BXpW
s5UMcgg3KQCHw0HSuUVbt9EAJAIfmoYEYo+bLUeDywSkWlAnI2afiTw48xq8X9kpjhPOvJHN33hm
3dqiPxCT2EXF2Ri5skreC6lkaWRqdWgGgMvJCj3B5ju3ai6qeFcl4k8G8wk1r+2u/wGaLwtIC1w9
wvfWViDMmxtFOyifi9uIXGLUwN+0UKcGrYf39M1xPQ8wSg0HV/pW3DLW2pdzzLAPBX2537hGCVLN
la+eZ9MwgLhc3SqeTOLePKFc3HvmyulaSwmhmvl2owOYS5n1OUr3MmKTVzyHSKTao5ZsM+MAgI4h
a2g7zhkdq+eyso5sCSCB9uWXii5RWGL9T3FCRONhkqnxOyj4A8zg/JvnMkt4XoywFjXYrpSpjXzs
L2DDbLflChZdD9hNq2CuzpPStSFEGzs2706Z0DgwUBV6FNEDa7gib8bG3UfXTPvwPv22T1MHT4hQ
ZLphZgCsaoRa7cxj1r0ifKtLeNL4uW1koNypJd0ff2rnaZTfZv/QhJLi9ePlqpB5YK1YebjD02AS
mYUfxr4sfM6ql6yGy8LnwHSbX9ZWGZ5OrwWI1g+oovcvreEUPcW9bI8tDT+1Y2b6h2WPCkYWwW4B
QXDBx4pEk5FlwhySuGxCwLsItf3V9l/7CDSCdVQ5UlAKF/Helc23oH2rV6x5kij4iP3eeev83FvI
jj8gMQsjJujaSnSSJikeUF8013YfncgdcDhfDtHxQFOaurUeCU7ULFA7+nvMxWJWdTh1za+pemQM
d+cpaNePWu80thvWhfNzmoYpeuYFGglNN9Dxbk99V9lrr2Ek51tE8VD90lUxe1FIJdOQEXHZuDXt
dkncwmu21Fw5b/ZmnY4e/ugidzAQuWerG7x7uMzaaeqJaHpDOshqKM+WRtvljK86RSiLwdObELFS
LEIbxkCFQ48ojvWR5ZUV8ZrrO/8gu5jhe/RLJ11kMvxpM9X2MFvB2qSttzVRqW4jaarQRFNfC8wz
XwrtDjM2sqPD02+aC3qkOcjaexv7wCVY3FGEeAbwA4aqsFxGJbuLv8LWPMjLrnJLdHFiDiDnBxyZ
Tbl3yBrCkHR863EkKMsZg2CBbUuHcHCqWFnRIZVg+nwDN2Y2+KW1FMEc/GdvT8usnvV2pZ7BiaTp
/9UUfU6TEkXZQ5tyoXV+Kmo6KS4brB77GUTtFw3l/zWlHMRHT7xBRiKA3g2YsmrbcEiTCaItNriS
t69HCXlwHe9ufOcdWuZQs6WfzmqFrMRMnQJI0rzc08IIsdBdmnkjDLJYokdrVdwAA+qBRZOmup6b
xQoLKf0dKKmRw5cuRahgcYgHEW8eLAAUE0UlUxxkfLXSmLjNhNM9+chLh32gf78f4KLBKkZP51Be
ozG2x2HAJZRwwnCHWNtjmAgC9MNkhBOYHVte5mtmqqtlO83YHv4r52m4+I/7ylw7BiKu2Jphfnj6
2Bb3xokq0OadxfR+RtOSad5mAbYHlOM/yrFryzXq9rdBRFN8EkkpniR91ouP8prl1q8yAXxGfXtF
OiBxw9litNp6ZprPfwmxxH1JM2OYqXkTCYGSLRQyJauISbOWsfi1mp2wkEQP1jLMgpmsgZ1X21eY
Sovv4bxPWJVQNMHOLr4MBzAYYsk6i4F/UhEkJRVNZoX1ROVc/ZFlhsjcL+esiAyu2Os9HKuheuBe
ZB5oC7IMejjY1vg2iLEEdZd+JZg33jkLO2r7RxzmAqNzCzIYKpdon3JmxsD67Nw4pNt8Guuz0BQG
ERNf/e0SxMxSYhpz5Lv8shPupbb4b5RY0vePLceni9XVo9X00Fri12h1L9v1Q8gFF/bcQCWuXU+H
vHrxjDNV8vejpwyZLJHeSGJH2W8zQDSdzpu+DOA/bbQ558yBzmLSeRi7kdERAGeqHftumL62ANvP
yMYzyb9nAKFaRfYsy2k52ZbWlsRp0Oj73tNq1EFzHBfVcKhhsF02Lx+oXo0vBna9Lby0RPma6ILG
5aqfYpCsWXGL5izRnvBRv7z5sVLSxzlU0HzBLeUuQpJu1vDrAzaYdgysdpb4pf/LC+TsVHfSVEFV
mkZR7yy26pGyWfQJgqUV0d8sQUPqOpJHY0O7ri5A6ZiljtgUJ6CGfOHdDS6jw41QPu6zZO1ecLdm
SmurI1tQhgDfLgab/TGcaFUFUxAaX8F9Otcqv/0k2OMyOd272AVtotrwa1vmuSMOOUeOlA6YGG7o
8K+0r+hVdzu1TvSagpyTAydkOHCU6pVHnKXQxDQ7RiQyszmMGZFJgfQ9YH8JmlhFvX+Ww+95Icv3
wvrhkhRM2Hr4JLNGkkw18/pB9kNthj2x+GoahCtBJ4li2YFgS3+X4vRYJ18r6+wFc/k6/7mOnMFL
mxH0v/Af0nybigNgrej+hhw4eiehW0C200WwV6SvlAot3Sqio3kqftCXh4uCd0ekIlIUrhi7t5Oi
ygFecIzyIFYo9O4IOOHWiC/Fe7HG8jiO4/B5Dl0BIjz7i56fAULzBz28ntgqmpoSBJ2pCPE4WSoT
FzOenb3uwhXEVTCt/cBLvQu0aVY5DEZ1AKZuZKwxs8UtweXvldbOEZmcX7OnLhBBOsnyZDxQYSHy
NXDTnYOmBxOUm+UIlGH8v09VOi1q8nh3EG2axZ3eWlpZgCOLwd6hso8rZrrwE5IkfTM3rJTTCwhL
OaSmizoGvARq/QZiUXhdlm10L08BkMYYmsU/Oly5dR3727ViS0ZdidQ9NJV44vCGsTQNRHYq4iLj
v7JFEcc/w9o4cYIYcW6R2tYtiqboCDfjV/nGUBzIyM8dhDR44wXpcBHpKM58yEgCn/tI5quyBynT
E7cSnWc+UWxKezjsjIXnj9idEH0uSsDcRe7WkCykDrs4ZZJ+Zzmc/HyNdgbRQjabXhqVzplkeAHK
Q+dv7lswfnbclBrIHgoOTssOfxCVjXMqiTpr5X0g3T8r93kqRuP/Brj7BCTaAFfOWBxkkzjlftiy
8OECeqU3/XAGz4jRuq0g0kskw1ndHVjVm+WZQboa0mgjUyzxqhU0PSeP6b0oEJQ/vNWk4NgOBBc2
gw2riri7or5GjycQ/WvhW6oXkm0Xeqli3fZsEG21y6lArsUTfgG3Hz+UBVmxR4RXQttdBwPnOm1F
yQQuyqyyYGShY8lh4zg1Fac4UdnbtreiWC4XJh6yz5MndxZpqyu3tnmJ8vUcjhoUJ0Qvy95L4wgt
iIpc2LPzKYIKyLbSX/n8P8VmjoernRgbtefrUvGxQmz69skVT88W5Z/PRMI607xyl/aI9ReoDA11
WPytj/HyizRiOS7dk1lC7hNnwCYsj58zG8TFjC3xdJmEOfDb6KEheDO3G7hGdwSU0zCMZTmlSIm3
uD2tVGxqUhBlIN+46wTfrDN/X98MfKM/8Bpn9Hbr6BiQNVElCFpn6FEqXWaY+peXxZhJp63Hq8JH
J+JnHiVhhPI1BP6RfGkUbTW035Mq5egVzj/+JbFWdn9g5Z+Cj7Dx/69l+KPjpvTotIWXXwjH+49D
CNUKu3r3nIr+g+7LOc57LykYIpab0O8ctTezdxCgxulOaXSI8fHmNgiMc4gfNyK4vKoQqy2a07Yy
hn03/coWtwyKignNvyqgFIwC7+N6y3AJxsRgUqRiNxNvHx1EceK/PFY2pLFme1pjyu67MYs+mbZi
dSf+/Pk9nUuXNsPCeR8yBu4umq0MSl+Ijx/x4pEkuc24PCWBuYKMNhx43/RY8anesg79Pg5JfAei
0pQPiweWla2g+DX6Dlp0cNFhBzLlVZTXhgSyRkb7P1izsQ2bKznB9n+9gSUkvWh6JrYDhjxol5mf
1XNRxSm2ly/Fysc5z5UdSV+DJ/H7helCssyB45c4M1IZRxWD4MbPEomaYpe0KKGd8YjAqeQuJZAu
GdTEQZBJQm8GkSxffYUsmkPXV2AuWOy4r0XV/avoaK/31bwy+8hEnyjpdbvTxXehZs+bApN0uq7J
uVtqUYMgkKG1NlTw1DaS2X0qmIWKuxWJSOSaN6QUfobdUflRkED0MtvEeXgByfGlolWDiooRyWNT
Tiae9imcF3ac/9q/uFICmxCaZuraqiMTcyI9bPMYo0OEEEUZHAeW0bTqi0d3gTEaeHqb+qleWOmS
7gwFVItOiRqhbXeMR+Z1QTQtVUYJMfeBlfkIc1eYrFuPPkO0PSbbd4k3tBCst+PL4498jEpsBx85
VS1maibUlE1Z75Mf224l+ODJ1SP5aJYzeDMR2BQwrwNBvNFlifSMVEp/gucheh3XRn/e3rnxnjOY
zwin9CB/aedT5gxqgw11hXgAfNun7oRCCXwxMaEnIQ1onYCE3t/S1ROK1debIm26t17Mc9G7BOR/
zEgloDy8Hn/zu6sTwY3usmRfaKyJQxE8rT3s/gD00EdQnYYPj1mDY8iDwq/lJ7lqoiUOHL2RvNMD
NPCJ8eggKxNpOW7cKqfBx0ttqdTHkNfJ4VRI/HtPRfC5CnDNRU1ZzI7dWi7tFWBxKSMekjVFb9XX
tpAP9acjx2QM1j7DPIZfcpHka3le8KXCI7SBx42Z7SWScVuWyuBwlfpXZZh5UzK7llnK4ELxEr/k
K1Dkbuu/q5fKjWdbn41eHiWOfjKFoYEFwvNXiZAKhkKHt2ofQ6wuMEujWmubGpVMYWfGr03vMKZ5
BKHmw2BV0lKYEsnXxQUNQhqgXtSFB0pb7HffCroCinCFQ163HsungssMjfNF8JCkf+UhggaMOHtI
Gz37Ie/x5kVYbr4/sDco4ADy/qKXXbwuAk5IbOi73VbjaXbrWab8+tVms+6npgo9P9abhO/rXxML
wX1wQZOTcrqOnn3sZFRLALwlwPVMHi72EGb/dZuIDQDye1HhjWEgi73xqHUmZOjILrORA+Fqx779
IrUXtAZNZy1gdEw60Wre+jzUTQJHEJ2ZlS6gMr96ulYfmdhhXdzJyWVSCUoquLDUYEnspAf3yWQ1
O2BRj0pJfMkEywEvyDiJY7+It0UPVblgB9Yo425CdreVD40+sBd2Wb7WuwJ9KaVqKX4RvH1SoNb5
7r6xkZ3SNRAoICfLbWkWlh6UgurRxn+2+kM3smOmBhz2DxNLzBlT90TF8eXFf10gECiLCgkMsIpi
s7THFU/Z1WzhTorK0g4IpnPIn6Vsajf2EtD6EGlyeJLN2jbQKyppiZ9fjBwKDTUY45eJYJzbpDRa
t0DoQh6LrTyExhEJrhsIBt/pW0ZsexiAC9idhqbHI1Fyd7zngGJ1vYmSDDchMgqjlMPYVQTmlAgt
DdOMw8tFNiah9nWpkH6zogWMAvyYCBoBp9HxPA2QwTwoDjN3eBH2C0dMrdb46OPtOBzSJroADq/M
1T3QZNnBdpgM8Nl5K9XHPtKZZxtxhTbuIRaiYPXKnrLNKoo5qEmG5iCM2NoH5LHmqV1O3x8YPfUG
FL0NJws56DWPf/se7Vqj4klAvdsH8l6C65fRDYpd7iPH8Fl3RMMyzoDOKYTQa1FWyXxxFdR7OZU/
6o2SfjehB4+JNEuZzeQcwEDU2z2pIT2BrtolauyFJEApysPIbtOpesQXcJpANg168iK/t+XnGlYK
Qt6pty0bB7lt4M+47Kt/W0chrWUGJiBvQsERHG15iKItsJW8nH++4LglQ6Hild4u5zPebsOIK2nH
Dy6NqCr6hBIDrhgGo8zFnNZ2T8SaNemgeKgLchzedMk1LXmIo/xP4gtBy8dFW0ZYSNbb5ICJ1uWj
NuKp6pFGeTyjjB8BdBrEDLiUfHsJiiHPDF879Q1jTECzPuYlBYyLj0+llqSVe/+zbUrw5Lzz98kq
Xj86MhmrGnNBsINclk1XUJ/fl3Siu8PrdqUZdbd6LnjxtYMqIVXizbSLi5DZBJD4DXRpFNJBsfy7
ZTYQZgF2VGw3J9HIW8BmPv5GHxnmUjJn1cYsFr3VCYMF42nsEopyr6RMm1ZMHz5tvISzCHp0NRda
bj7EGJlxzAW/k9q4pXpGVaXFMZJ2SpxsnBP+XBTufyJcW4UIZB/+dkAXJrHRheUUsUU0WwxhipxS
OZGKUoYCSJIGDXS361GGtINifU4Ck1h4wuXSfoGhOAEWMCbwq+fLZ0DF8MN0HZ4j7+5p6h3U3r+5
ne/3Me6HXCj6fZ97B9V0Iz6XbYZwUNM2oPn4Bprpbj0bNkU6Kh/Je+hpn3/jRX4bAYJuTJQmtfh7
g6RH04vrfESBUvdsm8GtEDuyHelJp+uZ2N2JMlR6Uc72+KdNhlrFX+hwi8jM+i9hy6H0kkA7myT+
evlqu1BajMolzrbaWnx3N4xO0scQ6/GppDV0RZpS00k+SCkeF4cWWzmCpjlsxDN7lJcWh4i5KNPz
icm3zvV8wYzkJA63T83tdwPu4HGmN0qOWNXCO+ziTg9janKTiCRTF4MGHjdpiymPTzXNDi97qQ0f
6R19iCyLLyLP7N0lS8Od4zHk1RJ+hVrQlAmGnhvL3kYYgpj70JSHbzCpz0zUu6oUwDeTbYQgwO3m
qhCFlXiwqMCVLhvFqlYtDHM4DYp7Oc4Ib74Tyfj3BIa8AbbolL58xp6mcmiGgt4Se1t9YB/YZx42
paH0qJWmaPbL7jOR71yoOlaeCrLftElvkCs5/tiLFFGBcaZ03tddgyoORJWZ4Mg/L4AeFjwBMwP6
IYr2HFzqzgnpxsuKw9VieLFAMazww3CpmYlC+QfoPfZcBlcxaLz3R80XB43fu38fxSu//ltp1QaI
0rWjOxZenrEfp+3NlVrmuKJWLvX1Ku2DwUTArOVCBfngKrxss6uvqPwObNr5U2I2HwuOQvvBBXus
SUBE7qWq8Dkb/jFZEhtYLNMvBgQD9UU5E0T4G9fFcrf9kjRNCRoSdQke/vfce85DPa9WIKZTW4KZ
mZZQJnkUBDnP2CmDSvgE0Lyve+vtL2Qll2tT+Sl1/otte+M4llPG1/Zz9+zC+UXt+5O8+W2lBFjR
ehkvsuCbgZKDM/lXZi7+g+PXAmJpolBrwanfTbccUmL0b0tVqE5ZEYR5ebIN1lNH/wDBo5TiMEZZ
Tdgk1RbPN2DIXviEBa/0tKIJQw7vDOHUDmo7fPZBxv9KTTNxrOIAzeCtk3LOrgBpoNXnGTHpYkxH
C8nl3iTg7TVX80qD4tRF/+vjr43YB2So7PiO1zghlGJ3HmmjBPDNXQZU2OoLAWA1TQbGUsU6adGI
KIEMZjGXGJ1gKyMz18IzFikefBXnRH4sD8Htv0db4mw2VN1CjT2SnpUnjxMlznzgoYK+R33O2o2D
QPJE/S2GJLnA3UlmCVuMCK7J760vUjhqwJg+39k4F7st7+HNuvd914FYCzcUJJzwte53WcgR/IWW
PJuxv/QHXb/9DiEvV94dUeQzHawnFhzXrznIP/RMretn1jdgt9ZzyUFC90m5Gsvpp1YHHnRw5yxF
mSHs1QTS2XnqJg4p6NtVmBpJ8m+Bv+9AkL1aAs7QHbZYPlhb/eQDGa++8hd4/cVCX5zCf2dHk1X/
ufAEFvYLSrx6syNHpPpAaqg96fEjiEHdRI1P8qV8eup2Toif4wxP6c92T6RP/B261KFbVB2kdfPN
uaptbvP4qaomz3Es6kvGUhXs6X39PFTL2Z7CUuAng+3CT9KJfJB+CY/xLFVPtWr4dhbcTEZ+k8CJ
+NTbg46M1cFbHUeu1WKULVWFmLx4Jc+me/PySvrmJymFAa6y8ZHJgAv7uMk0hYevXuOD5ivpf+XP
8us2qH7Es41iMs9And+8YsL6PloW39WVdPLf8SzAQvtXxE67Cfew8xzRcykkix0XLNpW4oXB12Cn
kcVls8vSwfwxmV8LYYQvmXzIpA7uRwF5Cp9sSfmTaV4DdsyAgocaTV22QqQDmvIghi9CH2Y0vxRH
zxnzCZoLyZi8Kj9LbaGCE9F9kBI2SrH6GFmJ+mA1j4FhrUqQUom6Pc0Hl0H+ZV7x+XmTkWviGr+A
ab/CRKbwjtGYCm6e2F1c+dze4SUWOz1VKAy35dh5IsFpVGQVlYkCACe6bZEi3Xe4qcf+jOLjWYDB
U0f1Su4ppAn5R3uXKmri9ib/eHs8VcRKvBr7nXgsOWeodSxZF2B4e3lBx6upQom6qES91paQYgh0
PjWIU6GA5zo7Uoc4sCg+i995tn3zBUfY2bPF1i6cFAF0Fw7DC7dRUpOHVXrtrAjc4kUOmC107S1u
eiMT1rPtqcYazPS3BxjhRC2aV09bIgOmpyfaJOQ6JE21tG3HpimMl1l4qk/WbeMlM8z2BXZKq9sY
kg9IpoD5rW/cEfm5x1Ir8cUdYikYuXvKK0LxJhIPBncwFsY1FNxMgxTh+JFOGOdDqEM3AhEdgI1s
gpcFWGi087Dhu0Jy2x3z6N1ZO8MHiQM/h0TuZcYcyDymHxLry57v8rqXh17gFpXJ4rdSxN/BgfjG
1xkVMk50kmuc7MQWtkPQtnW0TUczgZpF9o2Zk7/MLPExLQ3XEYw4fOMo1ebbiyJMBq3b8Z6XVtoh
nIT4BtOA2f+/xYDASQYxwFqd1B9LUhzIe7SDK/xqqdBKiAmElzO25mD9TUHMt/EnO5hRdndfr7LF
qKJ2oejxrnCKlYTOP6rDnHSt1WZs0V8AtYZnzBD7krVKzim/72Nnm8jVYU0C6vHTt/biqmj7M14C
60VJF8k3sH1fV3kCZBIC/RVq9uyarbSMdnEJGFf9VuqiiziUAELI+irFfwEalcUkt4xFnBstpRDm
OZ0tEQyHa9LIG3pMH6qtqEiKy3iU4aVs1+AM3pzfvZrB1Bl611/629P3C/rJMfUl8EPsEktLdRzs
RTXm8bhvzqiRweO7rf+u3ZlKku7CQNfN9x1FKGbHs/jNCusnv9E4lb4TrXgwm8WuOLi6oOjjSXI9
XTQHVjDzVb0RX2RFPVKKwwFIqA4UWJbAR4mqbNt4q0IOvDUN1/IhsrtpBMWqNOshC3yYm5k44Ke5
5UQVECBs3hMKcvl7h7Go6/i4Hu3AVOMeriw/gnxJSRD7d92sesMF9AzMe2MstOqh7JPLFZPR1lDJ
uvZW+Eat5rtBMnmmZCdRSQsn1Y4+bXKAnrbCiU1l2YSQXyb2TbVTUKL4grWgyJGaYeP7LLwCc9Wg
4HFad2AU27kOHMM7tTq4W2HBI9yt8Z1AbFpmK0IwjdVaNqGvlj0Ns4pwL1+vnfmosYk/inpl5Son
DfeK5r93JrxA4F9DwCnF8Trua9AjeRb3XJcq5m9diuTXHpPhIj/9cyPBGlOsNLfPyHJrqoZ1mAEj
yQrZ0Kl194ELtlAEALs0p+RXwURLSrzZZlOgSSz2avE+QPn6TS7G4idSkqLoeZqlvLbUugekLUgv
QX1g8UYr7Ra0lL6UBO22Pg8a1tmljFIzWFEJMdR7/NqOy+eF2AKWBulugWUXb6gHy2/lDIDWLJRz
6/0p1DF3qZ0iiIVc6k1BXBLiM55M2jR93TCr69A2T95jO9+eKJATqxc0cU46Qp6wotPkkq/FZOcn
z3d3Zp+5GspcmhyA2OeuG+97YB9dcmcUHHkSIf1eShENe6wyIcjnuJGeWNssB+Hhy1RD7fBXA9Cn
5uXaTJ8FDqMVgwZ91WTbFsi6EcfsGdGSz1BkbMAs2bhncd+bH0CtnF79d8OOE2ZRdolIF4I+7lT/
id9m8/KD+idNCCRwyvv4g4OxpeckSV1B1CoapQr4JLg6YcR+DdTCnuj9U73ELTrmbvXa0tkBZCgu
eVQPP1KgW5lUiSug/SmO9mHlsx1eupUIUtAJZooO31N1lLxnautZl3/dcAuus/TBAapQlD8S5hh9
hYdUPUvbVex9qrhvrYdzSeFJdcshlXLjMljB2gemLA523iuqarCd5W7TuDbd8mMAvUzpJO4mPSxD
88z1Fdksvkesu9RwkU92wQL5xgmkwYiqajzRDjvCOcPY3BtdF8Wxax7NuKiVYuAKfO92tv6CPhms
z9pkQoN0FnqGEDAavyas0BzCvUF/80ylm2muRIARmqVxkPFFM/sy/YjX3Lj2HUxit/CVaA4iYkbg
4qtCyj8+iCiNXAuLK1TRwyS3MHLAwsK8EzNSG9fCN71Lk8YL1JOfasD9I5WqaJblBwRBiyudhatT
+tlCVvRvtULqWxo6GmQ6gOs8NIecRKHUSn2t9m944j9/E3/juetdNKue66dts1lEwtdhiJ1jNnI4
XznHme0UQOPdiNzfpGEosbos/v0fu3UgNEdYUKUSbJJrjo0mgLwszMP61ZL8t6p/EdE9/wfQ5k0B
90quZXRH62yIeljbW0FpeYiaptuZZKI1BSK0mxDm8Hu536I9755+bFxEIkTbCM5jVeaP0zF/xF5X
i35Eo8aBaCD9vMYyBEeIiR/ULBXvbUou1A02fnNvr4g/+xtUOx0SLQ/C9GPNcPY9k5eXqYJC8jur
eSVVJ2fD36Ll6vTlpBFa2WrW5OlCPz5AUSeuUmhfe4AmkCEwK1eFCJjhMn5/ZjNxYz/9O1LAyjRo
6SFeO+5hEyBsUmcFhmkdZkHlszxgcEqwI83qHnMbw94iltwWxSangKpbzdH6llFTGDYXCsJxnLRf
4GrdAfQzD8f//PIrzVAhd1OAEeLyt2eyC1yYVkgZLuuGZDbBSAOKsBCxeqJXQhL8AL/V99U9BKxW
mxguoiJHgkAjNuW2yn8p6ax7KNmjVBz6E3SxMcvWuVcrvWUqoP4sUZrrqT0/7SfKIXcfhXPds0lk
iEvrMfalqhKJS8P2JHm3ts4Y0pfhgROpfn+0xo1nNFxVYL6ACKd3HVEegZGN/kz302VNlOXayf2c
b7/kwd1UtLDdTI6+AsQQurjj7QVdDRvipbDgbJUNMJ50o8Xk6Q4z9vBWd+OmbfHCQwHLdw+tr2qW
DVBR7XfXNXC4MBjhF+LwOcpPV1nBkF6fx5hvKx5Xw3MHSI31gRxfPGPzNQjnf+TT+93H/p5blGzp
SWzqN/9BtdYMupSV8bATc1QBK/vwwiyl6iZ4mHll6U6iWQEeohlS2jTqGpYEWhYWwVbOnkk77YGL
4MgbE9vWgXeHVWI9EzRrHgZBIG+YPHY+mUmOL87IuCqRHu+kzEduA9Jlw+AvjEDZ36UdrkwB1xRT
F/LyAticQihvRqnUQ172Hbrbn+op5jeJHXIXpCRhZ339ec3h9LOmQbkkV5jy1WRItjMgmkXcu8ey
fDfs5Wtq6nTPTqFnZ+Q4XkFg+oHMIPOEkQE3v2eqyKMFJOXHN+1MpLL3wAqGrhn3Lm4GriDvR0bU
rrq56K83S6jxaglzFuadbyP0R2tXMVdP+lHGDSz8Tl85lwTDuk0CX7aMYe/H0KIEX//99XaPDyIO
1NzHtAABsLZBFoRynttsphT9mY6ZstwzY+HhXAjeyC8P33FnYcqKNVHjWgljusJ8MOdzWyVemKAh
XxdT/ZrGPv2bRL2TfJFvxg62TAyzuvB0h7heEUv/Zs0yoVG8C+WSgwbQpADMt3MU6vpAMgkwUB8D
RgH9nfQMvfauLdI8N5r5xNTDXlUFiFVgfGE2V18Ts0dBhuMOjVu/Dw6uOGzP03LRITOIzWXJ4BFH
UWHhC4uONh2Oi9WdiTvJQc67BrYMDD+pbcASHsnDZE2qMOJCVIm5YAvNV19dfrVich2Qe5AxUOp4
imP2VBgUmbkPjx2UcDTMUGRaKoSvghtLqoDf3wEBxNn6OuwzUMLOiArmDR8yxPque46YtYAtfY0w
Qhy+7EE8osKubvMLdmLNQ6zN1fxMj41usEQ1jNTtwLw0qfW18NIyQGg98M2ktiYehypSYLefTrey
+OuuG48TKtMM3FzUaRe5ihdG5oEhppGs5+LWy8MyDNq1VMXvGINKoGF28JmfbQrsIyBiahaM+e9k
oADWMXNKn3ofGTp0jR3Ba4xpaz/pNDoW0KbYgDjvFUXsiQb4ZN/FFxxwIPuEeoIXOTuBb6VVQ7yJ
nxQUW9VUqmmV7wBqCM6axOBK+Byxp5pZPxQ25Gg8w2Ipc/aw2PFPPzlvbTgJeivGOAHsv6H7ZTXN
Fs9K58aA5uANn+fy/YAR9m22BIeNVkk0uztEygGcmRNrwLyaRdE5gJ4mdgmWMs6CnVtpRaAPnDC9
qTlZNDJ3UtU4jYXCDIK29Mu3Kki1AzshAJvvxJD4dtAImvJP8gcD5zKXGcH6f5zPdTQGTMhaFiKg
Owo2YoCPfBrM8fsN6dfzqmccObYC4JQogRHM+3RWXePdxhgld0Uxxb34fawBtcUfqAR6rvgWB2GF
3K3yH+iMiUuWV4JosyMEj4EOmHzRYZYnB9uLimouutypIe6T6UXGFSMS+KhGphJbi6S+ojWkQh57
AGG10WdAYi6XQJB7xWUoXIygKx4I3FW+2UpHVRspDioD9xYsb2LtcdSPAVM9/bx2hhNM4HQXGVWr
VifiF/8CmwX7dckF1929oxMQSyYlc0k1Fd/WwxPYSurDYfahHpq93wKj2aUUacM3inPDAjhenfcr
Ng+DS2CspEQUyQUvVrNMVgQ1e9qcPBu3xuOC+vBIUqxjzRlMr+6IVzGoQH64AJ45mmKwJZJ6ZR41
SwOpMY8swLPQfxZvrgSYRpbJ19UAU9Ph5OdfW9A9FIb1jJSWhjFSpe5ylhqoupmrkcjpd7yFSZIG
rFLwpOdnSIPx7+RVZSLVQyM9UgQnQ63Bi/MxSAgV5gB5NbRCl8M4RoT4jMqOBh0uP1vVxzCdBwqn
gL6Rp473aVnjJKE+0XGanf6NOVWKAwGiroHx0s6s0Hw3LS0uC2lvgiw5iUlcmEmNDT63h0jhw06N
Zsh3jWrdSoT19qcVVUfi7kucnz05XVvu/4tl1L/BehibexNLsjtxuD2EZbRXBicMxcurEFnz6SB4
LA3s/VNxCkq4l6hAd1hl+jCUmnLexH1AvcFKSGv+rRNdCGklbEH7mOFH9F3WdYjPlcFI6E5kRGFu
XsOwLLAn/dKMVioQCUhJ3Nt1+FWubftRy9cGt21Yj+0xpehoy09i1Duwpcux/BKoPjHjeTrEPdIC
U3R5EkTY7Jjw77S1N6xN2trUrdYRyzDtBuFCYT8gtpGHH51UQ8J5L84Jk1Quzu6JlfDhpu+eoyR8
Br9iI+2B4/+QearBMmEpHiNiSmhlaWjTGVfljXe1dyd3DNpXPINsk8YUKshFIz/gU8Wu2kA8VQ22
sPXwUyrOc1WbIAQKRePc9I4PL2GymB5F2c03M5HqTnP99CNaYq1WbtS/81jYbMdR3goerZmWpJ76
0CsGFkHDXFQWpi6DhVBciz+HM6/pQglqD7UOAxPFfHNKH/TAjONXQQWnjLLKqW3xN5Z8PojOYkQn
h1XXVOa72qhu6+/Kyuk4KB2weptrfzCrEiPLUIvAdp1h39zI6keBVHmBUCZCZWaol0RiymiLUe2Y
k/Ae6Ps+CvOg/i1X+biIvvBoV25ZaIOXz2TIl46P/1B5aRh+pL3ilnz7mKq8GLOj3KllwINwM7Y4
d1goTIMeX9MqESyyrudFqHqclNTOlME01CykjIQvxh05orlv2NEyLfpw+pJH9jKaOjHDjEcc/30c
IlXBmlLj5Y8oC1403mZj5Wo3g/hDudmOaA+otlub+p6mohOXUCTh+4khWWU2IrK0kKvaXkEAfcIt
LvKSr1ha9MDcGQ5sJGxiaUbm/r/3Brak0UPEPtzwkNdy7HFWFh271QABq4R6zVHdPu9YdNEZq8a9
YnTjGdCwSM6lsFCJHsT37sbzwhsq86LUqNkdOLjeYmd1fFd/aypvCvKRYtS9Fp5PNaqg8V8FJyr3
dvI3PtS+bl5FoastbOSa1VKZL6NsLGwU3e6vlZKqMRo+1UYlouWzyaz9dBZPRvdc4C6he+rTyCk0
K5+9j2oUVmecOQm0VTGRECvXUYIL33cxuTVw0KBUbvizJ9jWeGnWmE0JGwanGK0CC+XPnbPol3JQ
BVlF0t6uqTVbid+6kBSJJVtt1Yy/CYDt5uK4gkGfIECL+uiImQE5zB3c4dvjAZbd/44jBx+SCApB
5psZsCMuxpqBvhO1Jx+9Fl4YFYR+8r0SHjq2NnLR6yeevvY3GLxuNQdVwRXj2WeDmNGWXMGTEtFC
UJ0+FqD4S5m3oE2Gys6yupW67XISFttJKP2lZeU7pSjsBhuDtIWkxyx/ArwVOw0UoU1nQ2xmEXJK
hMLcC5hRVUu3zsRzrnQ6HNDhOKM1es9mLIQeozY4QZyPppsp+vKWfQaRjQlfpgyHoocipZq5+jey
V4w6SJJZcp1J3ClB2hKFL0Fl8e7jjFn0dT5ZktLbAaA2TMsyTDWd4oOWiegFj9yjdntikCSXvQdQ
+sCJfBzPQgfL8DxY6otaJep4fLq5xGcfJTSvXNkXXxgZ4bibKmnwQ1c3q3uDIQDQvZhUI/y3n1UR
5mK/YWKvc5uODMlQaB85Cks9KXrNwZ/b99dWQzhdc9KcnPZWzYtFkAFHs659SeNGRCJrPoCBcjfv
vBFKMp9ZvoV1vGcNePWRauOSEN7er4MZze1GHDD7U1OevyTVrNWQe3o4XHSzRzF+ZNG0yZtjTe1P
4jVC+I22dyPTOs36xTbtFhE41Zqy2QfP7NZMZq440MaXgXZpKqzeQ4+7mapGFZ84rz6W8eFUST1x
7DQ/JZTv9loQgp7MFqgC2dqIKkahpYChRlE0UeEJ71vAR5LLOiL9TIIJynlI8klNFpzngMoR48dm
cil8lZX/oehcWE3blVbHObkx/8oP6o+kunfYPnKam2x/LpbRg5iBjPgHxJ0WuTTqVF2hfTUcP3Ix
GROyHKVlEo+q8D8q1LGk+lV9sWGcw+V/gjSL3tWRUHFQA4My1bNEJWVpCxfxXFgkb593uNge938h
Ev7kJaTZcvcuke8eAfygXOfc6/EYOb4h9wkkM1qO62eTsQffnuksJ6CWuXDeXVPvhq/5C0GTwWie
qElkP2MOZg4yCmUOy1cmAboSmNLhF2jxHYRaF4NKibaywspzbm3mmqDx1tcGErYB+FtRJKqmAoFM
Myi006MlBC+yakbeI5ECLTYUYzJvdYX+fFOXm0V/Na0OuihPPW5rlspzyuf+O5IjOZ3el/5l4v8L
zEzsPbE71PmaNrl3q4SYhMuDVLFDWH0rO1Sl73B432THPoc+uYnfTJqEW1M96Smm/rvRCvmerHk9
ocZRLFDzxIdz6Hi6AsJZxlyFccAPt8c3v9HatAGvHdvpU+IDlgEni8a49T5PH79JxZ0oxqzQVeHb
BDY3xo3cqDTbkOkp2xfBHCxkofcPVW7a/kSMK6ZUfpMzl4m/Qr9khZfjHzNYjn5THraTxqdMgZzF
Chq6oGpuhW3nAgpMHf1xSXyS0ZQwKPirlD0ZwomZ2xDjicDv0AtQtmSOgdruUlLUhptwHnyN6f9w
dLHv79eq20nq9oIGkfaIspArAaHF+bqtloriKlQB626DNLBe1y+ERSVzihj5++rEb+VmbTpgTSBh
nzx+quV7LqOVIw5Xl2Gv4F6dOiatBCK5iGuJbQHtxn5DhUYTkoT1UFbqYP2kgg8lgkwgUgwqqkVg
6oL9xMrPVQFjE5d822kyPjX209qPECPmH+VWYXgL8zGUDL17chH5IzdDqyHVgIFGiE1Ax+c0YUvO
C0cLMhdVgJXP5mZWuadeNF+MDVSoCgIYyrhUmhLgaQbDNpiq3Zw5dWVVP7GYlhxy3JXtXhpS+CO2
kw9+Y05EzGM3exypmrlrFTqtXKHiZiilWw52zj70hS/VpCgh+bw83vQGzfG/Dgk2ThX+S6/Bbdfl
v+MLHIICpBM4c/tTcDEBtjkwYHKn4P0nNdsa5wEykOVlmsnh0Q+EHwNC7xYHxs4JYPzugT0oPHc3
2dGc9AEW7nrYwm+CZBu40B6Y/oh90u2TECqUx9yJEH7yNukyVBZHGqOCm6XTMZymRaOtRkOhT6Hl
w8XrbRFEwhnUKvtq4gWkW4aB+0eum0d/nxg220Jwh88De1LKO6lYIKq96MqxVS2e+9HGn3TMtoVc
YLbC41tyyNt2E0Y5d0ZT1RDzP+5IXd5++Bd4sAfJIgf339QyG7KJ5dI9l+gUW1BMKIGHGdbrnwlB
lstktBGwWp4ceDiwXaoZ5Ze6mH+cCdHOj9Jxu2UYYRLl6V1C1yXcaivaIHJUAntVulTTJf9ZL9qr
YuXEAz6UTl4EaUqPZctP9AWHy1bVPniCC1+M79jjbud1McABQnJvuOumShWRlMaJ+NK5QedPMlT9
W7JnDwN5oP6MiC1tQS6bwktls6kta7d5nPmc06Gqgjwvq25AUKBPauV5bL1i5caG+8O+HCMrW74A
xd/ARHMhbkdAkLYWBQelUQk37FkOs0e4XCPNP7D2r9W917tVjgzDXQ/UsiZEPdA1pm2kYFKw6qJS
DmRWrhZeSNqWd+HoMpSQeRzGYYM9LfP8BpqVLq8nQG2k8AlE5PIDMEw+ykkcUw6RhDgr9nn98MGL
Qkpdcm2/y78VIfVW49eWEYsd4hcARyJpd0OZc5uCQ9j7YJrJxG7feOGLn4qMsoGqHUUuQG9iOfem
7FA3MpY8kRvS6xGnqX5eCrzkmHoST3zyNzmmTkCXF9CNqQaw+esU4oLfjXFy/5HAbOOKoQVFrw7A
NQAkR1cxicvKr0r7UBnlvj/0ZuH2TF8N65om1GqA4IliTcFpM8C/PMFtrWBXUn/UYtkGSZwW/Zhu
85EPkadss8Y3lKoL1xkcnf9k5L2HKcVpTfgP0pLWxX/k8GxTKqXAY6sevfahQDnYIK0VfDEsK7qH
bH3qpS7GWRCJxIJCGKxV0guFxL8nTv6c/sJaC0QoaigbwOLESu6TGFvLuA61VKTkUewIis9cEagE
ZnbHcYJO7Hk4Nn9lu9oTcJK5FW6Zu/oPKg3R32LkhaRjT6o9VaGmgUiwpMkzbbn5iLVNs7byArUo
njFrpTX7oG1mfkxZijv+zJ2/uK142loYjEhkv5U/sZNIgNZISynOLIsi3sgaGDjQItUYQSIy8H/N
Rhv0AkjRd/b0O2KbprjMBa4qYVrMjWBjjCIrKU0ctSgwz6luxS6jOhfUkLzqxwXfzktEWLmTBomV
f1VHbskLOL5mSgUSE8cygsF+cJf8iGeEzMyHwtfMc+9RMb5m163wYyL4+SkfSu/ZYJ5RBuUE3SdF
Ux8Gb7tWL0guSPv1nSdIWsxMH/65fmpA7DtmL8h1g0oX0xsf750CTdfZJ2ha4mX7UFBYAbNcTCze
vsYxnuduePpjCD2uc3aMdxhPquYGUeQIypFUHCTq5yg9vfWsNjM2vZuTv3Ijag/7l5j/PXhHocaL
hO7zxogBWiRWJntz3zaDW6wBxUqb38pWh+Oj9K+rByfvkzEgzMD3nbSLhM5JEnXNzs31N6zxY4nI
iWQYFOKWIrvlJ2DCaA+7MkxYLM35EsvPBKJiel8sEu8e30Gg0ja59zfKlJyx3TduMtE1pa1s2Gx1
dGWUQ+DyS1dTPgAQTlY9padMZ0Jb1GM5LGb5LMke0yQWQF9na/NxEwZn0hUdmwzN4kBRb83+Pkuk
KBxHuCONt9urjEiWhQSXX+FGvnSYwjeWRhzAvwwtkM7ay4BqH8Xf6LZroeWMG62IAG9i7haGxD2d
fVneiMPmnRAXzl/mg2GiXsa+3t/9Cvorbd8b78J2K9p5Ac3IvLKq8dF6zZbNJ3lqBvMJbJ8DTp9l
ToB7nDXR6ld4W8R2C3n3XeO2OQgChXF88Oj5hdeufcmmQdqTPmgZbNboXYyqqC0a87au7UZt8sGP
3nPlgg0alXXJSjtfswEmydigCHD01gk4SAIjYs6DADuAdJshGrkm8l81nxCKAILZL/ZKuxN7wxrU
+/cpPqCFwpXs5S+IVR4C7jCOSVqC8aeL0afdHHHA/v6w5lpEWJKZeVUH+3+7IBB7iKKDdABWvjtf
AvWerxbVKuoCL/pDBaQXqFt6wSWJNBumJc0HVeU/mrgMZdh9C0tz4kNcFaI14HOuUtcKjPdKaWkS
of7o2I/0NAI6mL0QDgScEve7JLf3rUE+7wDUDCpCW1+1tzXTHw/delZmeQIQ/YxqvG46wkCpeETN
nODnYXyY3fawwn4bIOUc8BDKprPofviizgnAk3IUA78LVYOMMQuUMq8jiFf1MA43RhUdVq5XJ2my
0AuMSqGDIECBQu2VQCWgyULacuMWSKAtFxVYsLfA2bIVfm+fpMLRCST5fnbSNdbFvbAZhpwHhLq/
lIRpIQBBkzEkd2Yj+UNVnZONta/LKFZXF/qphx0/Q/+fBD/1F37rvn16qFs46X71yzUm/FVLaJKD
DMfepkvm56K52lyK2HAy6XFPAvheuZSXFO8+SG5wUctNxzhHbwFvYKsdor6dNX+nk0xOea618phC
7gg2+bWPnf2zBr8vPhn5U0PqZ+ODNUe+1w4bLQUdBs4mfFdOQeF9nL0mNcLNFJtg33B3upA/kg0N
7zLhDiuszKWt5FmF8h128P3fguw4RO4Br/WTCeUpMYvSkC2UWE+oYs1kxSi9iYWgoxFWyfB/YqLM
T/eYlo1WphdHs7jUDUpFn97p0mydxkLwq7b3sdUnKtlu6Q54oH4Ito4vgDzRyTx0bakyDN8SzhKB
RZU4fytoOtH/Kad0w3TFZjSBg1VWE5xE4czQ3fJdbSytHk4/E+hdZerqFK/H50OIZfoDc/5adDnS
fWhN8nEY0G7DZ0fX3tUnhrfOcUdsmrWJbttdAwSi7wXYQ46V7lf6o+qbS6wY8N+7jbrPwbBjiC3G
UaDLHNjhv4/M1S6FqHXYWEAHX8affCf9Wed0qTBCzOoOIPE7/GGCHCefhQLUMPnVWKgmUXN7D2VL
elOiI+fV2rX9BG6rebkKwcWDMblJnWRB6DAUTBw+Efspw1kKS9ldoSbT7SBWliGaaI/3qocxcjVe
kEDLSQi1Hva+EM/I0L5urC4AGddaaNEAEP5h5SL9q1n19+Sg6NaWrBpjjwNJ5PX4P3K/89IrZ/W8
K7gocpgPyPAGyQHZsAhGK2X13iyk0RTArcj6RyAlYYEOYhQ5AELWLhNvmgcZg66RjItltrRDMFJ6
IBQKj+4V4ALKMZwiEFaRg4BxRJnLqaE9t8JmXJFHYD6zPLs6lGCpnXlgcDX4TMKwugM/W4RWQPBU
iUbXVx5TAtTg44tSEoI44NGHvyxOoAoCuY9/LNDcgC5AZiS80MHwSYJcBOMFawTOJLDZgMzslTXI
2Knxwy67MbMR5KZcy5wuwwmOCg/RiKIJ6u5HQuB6V4KkeH+WARbOVTC8QV6fNSJyryu/GO2Jrjwa
5zSl0pasQp8Bg4zZKwqjCFHxTeN60kf1sbZaNirFVNnNk6GQjIMl6CtTJlRpxO1yFWRX8WfFq99+
I+nn54RXzV+tX+uHy+n5Mh0Qm6WZW6/ZBYJJM2HeQ+7UvDlPyunFKgH6JkFlK1AEykzOVeZvqVf0
d3+AO0BbnEEPcslbYJjDpdROgLNQCpMMjbDE1CU71t6H4/qpABqevh2VwcBqyO09Hf1nA2QAR5yx
4/RTtaGuBWo6yxI8ac8DhWs2Mz74D6Ei0amRHxVNunOxJlbvSZbaeTFV8BzbJ64Y6ReyZAtq9E+v
jeAVGzwrnbZ7qtpOikOQ1nYSjGGkXKFqUZCq/T6qjuCtbfCqopUlxAUlCoUm+tKVFXHg1XLMJF2m
6AFSrM7RuwN58vHpJ5DEVeXdjaHArPCSX9JTSpqAHOcQaOwS6RnQreZfVSH/voQ6AzqVLxotu76z
OIiDWGK2WeXSzUiZQVlqk4twAXfFROP0nL3VZmXWAeqXxAd6JYfBv0v2amXsSxfsv+qo9d4wOpx1
foPgGWWLHm3+ZPtCCOiNM9oFYEdEa+TUuOyhB7GU814LMZWNZUQzcCoNQfh/dlFk2aH3+RpQf9Qp
PRUM2sYvbmJ8/5qkCbCv8Aavru5jDH4+XCLevEChNKq2bNn9913BxwO8VYNDq22HH5lzDzO62YiW
KKJfDxsDyGJEV6Tg2p1GPrQYk6KDHaHTTBOm0SPKQehw0lV2ciLQYRvIhZeXAQ/4w5r+uLYTMfsi
y0wLRi06kCj9vHgFzLtezVSIBAl7V5Tn+9dMypVKk+AZ25FMcivcUT0nq+iwWLyxmpKyR1FkY+Pg
hTOGNm5rwzCOBpNCZp+wZhz69T36J8hpiJQmfYwNlkffsxQdu6wkdPBf5/ly1jAuYIF7nmxPLFm2
ZSm0/r3Pv1vh2JKRzDcwyaRoto0HVQxE+AaOunjjj1at94QxvAd6iSRieQh+J0Ck0ZDsNZkEabyg
Hlf3wJh8tZoM3c59hJEmYfoGnwK7DuvWlhqbhS/IJkCRrrd8QklRRyE7AAajCs5bJDZPBgomGgqQ
PEPMYDP0WjauFqVQFHslruKtEhyEiclskowKra/n4YJ4royLHLO8Eudtcv3mtlBd+plqTWioWYYh
YU0VATE3ZswWk6QaWd1S1fljLmgmRNRveiuFn4xCg4UCpHeX05Q5BVeGY9XLNYIeyIL11SxgWcvy
pjNRy8T7djzQvLa3ClTe0aXYBUByMvw5tJLmWnYVlkF1UuYmUjjv2Dk2tNUhYtY+ecd2v4xuhrLL
NL8vKNMvNv5m/DsncnfjkcBK9d5LT1bvtH9fgpTKSmlkiiX2mfHAFARz9qOgHDH/RXc+FAnoEsrM
lD6FIWQXzxpzhFH8ReVRMJ4OY40sBNKYK0R3gacfYidfZygvtMNLgxG8DZpyq60TKRXgmtxNQliV
n0yXYjA9u3jjnlqrL017wLHzqSpE/3qaKzg9jdLyF201v4gYTX3TgbsGc6HLowwTu1t+6DgNutLA
VJnHZhTEHy4W6ZjKaDeqXBUCw+uM/X+Dr9fjbpxrndFHrQrs5Bydi6wnp3s5/lHNmfge8BOsApJG
bmEweetj2Bin18X8ejIMuEd40T/WvmxAxYRs6C8l7ns8FdipjqhmXZIDpKNMuG1OzVVpMDm683Uq
jgcoiaA4wlA9T6bw+G7G4JuNsm3/cyFsKG6aac5KZIR1o5fr7e6wpE4Ef6iAib8eDPIMm0Ott4Bj
qRGaH8O2mRYu4mvj28m4t76jZjn7aDAD4ImvqqNrU+rSL7Fo25MYkeEv0477aM5aQVClyJi45s8Q
UF/YDJoC3DhSIzCJBommAns1PZTH/1BTE4QIMq1qtniyuivmw6rWKzekZiqVWAIq+D/+6cE9oVwn
vwiRX6CGnxB8umqjFOXOrOZp4886LFSCq5ftcE+D+J/cUalhE3KkqPErT5Y4OuebuTKSQv3ZKMP3
iM4ByLiJmH7/Gb6Mesc/MKcCJBe2KPfLt0Y5nbdcCfAA8RIiNvyDkBGmpFLe30cxB5ChvSqoYpJ5
gh3Zx3lG1IFpFYdmKo0Qkd6qeD4Yuj1Py0QApRfrmAEwNXBrGak1jNSTUDMnhF4wXMfKWaGs5dW0
A5GP+1JfAQ0crWEZwKIOJ+i493AxlqOLOe9SYVGSsPtGskLcQHjx+Ut4J/VB6aRJanyU17lDnB+q
vkwh7Y+zY9ePMjnLfsH8JkXQW48oUYKp4OCgFMnDsZ4l3xGPQhfKo3+uoK/UQTKBQv2nMu1nB3aM
5yjxMd93BUnsdzShWDob3dcUGOUzDzF+gg0XqKWScssvBxt91ESR3s1UA1pG6FLr/JS9KlyWPoRD
nAOUrN0x9r+BHpJGxhKVLchKRV2TcvmjZZc1wH7PCntt9fGnqE3b2+MUqcxLalUbgqQOCDW9si/M
EaOYXwZuwqhza5IN8GtYmTlkDCIlsTADX0w6+ZNVLxMwUg4pJBa2LtKYmLYOmibUb11tbTcojssF
v0Qmf86pBT0gqYQH971Mvbw+DZxjzKwufzJUX1PFsvNAhoz4K+XjgOYQvYBjHd7L5un2auOapiCr
Iy52Uinqp96OutWSS4by3sSYMYtVelGBY2YwEXK+SllsXmcZbPWAofMgH0HNzEpr0/2R0O/MwLa3
xraRwaq3uLmDIBfgeHbohfpPSVhpleWVRswXIIfBYUnKG+E66m7Y6cb4qDCBhaee6m+n/OWhD+BS
VpxnAxxMdt3lyofR2K6XQC/F7cO+CUcq/choblak9etcm8XTkpMHyb/ypRtV7knIebVrqqqRqzhH
s3R28lWBvX15SQMOEHAkiER4pR0tRY243h/Cqn5pk7NgfsfSGXbxtHy2vQKegsIxc/U/Joklvpcy
eWUB9Comc8RRshdPV1g5mLMLgenOqi3yMjYcDGtm91yATLXA9qU/riiJQ4MmFbigxPqK/oG/fkBa
0bJh1iJPIXAHdddBs2gHSMCnnpOzBVnfIWP2s1IEcAy8oNg6Z+6/L36s5dxSCvkT3v8c9ltoMBwd
iJLkR74KmGYJLKnu9k1c9mDdu1m2NLCDjmwCr89U6TnIqLTpnaIntbgkNoX6lpEgEGYPuDYqqq3C
YJKfkNvkCZF8YY6pVaxG3/yMeqiq8QGkQ+MCJ4I1FUTjK3tNh4nhNPG64PX4DEAYFMR6LsbIjpDq
/5AdDhO8YoH0xMJdIanhv07jl4t0J65KJYOi6FsX9rPgHS7GRk9R9sSrgBIpgSsQmhicFpZyi/2L
5n5Y3xcye5Sv6gUX2aiHwghSWnNuCy8GXyQu/1DxBpWhX7767NI9os2IfA7KQehRmaEDtZMF8aX8
IcvMFK7fJB+Hf0FS0Oau3UKbMyCFfcopjk0xbjUKWPHW7FaTXCRE7N0k6c6do3LcB8Xbgg3bWSjC
Jn6XH6Nv7f/kAXkQP0hJfpKfhy0aSuMzNN/Yn+wQr8LkrZbyuD2mda3eF3J4HmuxSVi3nDQGl75S
okLgANz9Atq0Ago07P0lIJvJp5TW7faSaKd6brUXY5+1MQ6YldYERWrZ694w2Z2SmpV7e/w0EuK0
jZI2XfUo0AgerlT6nscBNzT6m8pghMgiczcipT12xVZycjgZwqAxWoRvnTgxq90PRDiqMeEolhtQ
4LqMIP6j7UT1ZWdEPPjoDVU+xkNkGrjCU7zBtpVtTKUgTsK38H+vZ2L+NS2RuzOMrEEExIBy8USb
6D5OCV82VU5W7Y3XXmbnS7omFlRC4tEfBjve8GnNe2NKl3K7WDLPF7WXwLDEQW9CKwXab0XA5fLo
TE7vSfmWEI9PkuO5me7CtMdDHEM/5UM92S55RUYG+MeHGQ8HowBGoQfJYrHcVEyO2WSf8QQsDRtk
2KOFK5bIVnJhqzFa01ZRhKcAdFIQxTo1rV3BmK69RsQgqrNKrhomH5/yzmWCVkwmG9b3xcpRstj1
3shz4buryZYnSFOL3+9NrAIRVjKhQmElfEmAclGnxJoGk34pTYP0hABuxjaZNIRmW3mIgEfhdwRX
efN8pdgt1srAVizKcnwqaErz+hVC5c7CKkqhcr5HWdpSqE/dCw4MA9TaU6ETbTmlJxl4bmmxC3S1
sgOg9aLde6S3uEkE3+lffXkqyyviOv52IvTR6F7CV6wHndNpw1T/0p3CQopRCYbCwKsLnvX62GoM
Pk6e5ToHol/JFZ2G5MapMggW8JUBI1/zCqUCEENKrLfNrRHc8Rk++Vf9QWJ7lABSnWfydFvFkaQQ
hagur4C/VMWh1UebxeO+9brKr71muEElJX+n7cjYRvKW0jTHkC7kVFxSRC1d2+Ea1D41/ZNiA3Aa
Z7r8e4JLIrDKiBWD173LIvbuX1sxLGuzeNwiWjtmvIhvzwH9RJWZ8j+hvMsAqRkOmcrCeOWnmFy/
SFeM1/arR+VizfgXY6YVJZ6qm8JnaC/6mtw00Q8H1ofH2s0niX7uOSXOX0hSYxdEVEpckkyzWwPI
umwgLosp8eDMNJ7Q7rz6cBSV0zf7zJhCaLiejBVcOgIULx6Kak/EcHvTSXii28+jeoZrOp9XwVkO
EqfI0lJm/jznbtg4tvhzk2GMerhYF32tEvyeunq+lYn0DD1wITn/VaZkiTwdfoz2qCXFDeXU2oys
ojNorKZMVLiBGWs/kitzR15W4ZBYsyWEdwWRCNf1s8ff4u+4Tz1MnpDUCeujwfdhESqXTP+IP888
VFhoO2+LkNCFy4xfisBFXOAH/Usml5VhRGq9a7ULB8zVu1p45XDEYKtg3r7lpOgakLvm8yJ15QOC
5NACzGUcHiC6iUadjYQ0HR4RnGlXZuiFew5mcbFqmvG0HsdYYeRsreMMt4ZmKIR4cG9wNNIE+yU4
qQXvfK3MVYRVuCk7gXyhkFob1s7kB7DobXOcR0qCGxrQ0wP5xIH36gkHRmgEo5cZQylRpttrKFhR
MrJH1xo+6qRUYKi1EEJgdlqmXHZhfEJyb5BdWANJLFOTpRQ2g4+0XS52XdohXwc7VYZ963daIY4h
QR3iPd9qQHPdgp7iorV4AtiKlE2OfxHkUbh7xkxrEwKDmOQf6bT3xQQdR89L+x7LVWfKPLA6r821
SdPU2sGKqJUc1LbrKEQt6mbYd6zi9KhUD3Zh1kWi5f/WrcYS4jcr5uQqiePLoKhKVUAKhQ5QQj4U
aw2GQvnpwjhybnBm9evADcyTw7zfHLnDUPeuFg+DiC1jkdsJTt5GdqOhWJ8vy1QVUQklpYeSbj9q
ScxsTV6JXKQEf2kJtOrwZsCszO299J4xJDpAhxhNtCcX+eYfwhL4b1WVK3NBN05rS0EunfCBBrrO
PjQtZKPnY3+wkuQ+C5RoZkcIJZ+r2P2vdulypXFWIKZDbk9WQO5j05meovohg+2KMWZH4fH3tLoL
1B6R7iT/mxs3wqFdxEVt39CKLIrIbUAK7yj07pUM+2eqXFFkBs6B7D2wTzgUR4SRBhIEWnqJs8Rc
goQKye/tumGGIfG7lQPZKldfkcxZumTHriNyzM6YZq+WvydsEMiQkfsS8Pq5MLvtLQnO7Vn/SY33
T9/sUfwQpDsdIvEAbrlaQXv6hP0LgHfUd9XCArm4gLAoYM8fumZ+FgISMaLLAhgfOGIsSV5rjUXS
Z0YAgjFxWkcqfj84NyefRa8pNn6p5XEvL63m4MoxDnPPlrINenA/lo5H3B15OasSuOIx1TLmkJV/
RYjpTTolZ0E5A5aWXQAcOWHHb9y2OwxsMvGtWRfntQFLHc58MLacI86qo6VhFidoCmAKvA+0lh5d
3BvELQPjfIaSCzLXd2+6fFWPBBjeUQ8wckYbTJa8yXiX0VFBoIPTDvI6D0HaphwsyuyPcqMo5vKz
ljC168l+OwQNn/ReA1HHtAsNF3FzWFBfi61J7AVgW8b2ZLc6em3NSy8reTpnRlXk4bptVapD54Q+
QbWzu3MC8rlAlpBTG3l6wEzD5LbDFicW7n2HSL65/vIoEeztZcuGEOij2YcE+gpY1wSrxuO0Abcx
EkwZsV8N8ixM+7iyxtub+hq9zjfb/6yORzX+kRPr9YFrJ335iWpBqHU3Tcts7q/loHxnudgIaiSj
Xd26TlUMTyDQBX0fNC+Ei3oQsPyGlN/FhPISMfI3W+x0FbOFks5MYIOqDk+Cmd8cYxnfU0Nr3gNd
VVkOZtUGF4+iI+2YCAoO1ggkx36EFQbA/XEFPrJMhwiLGjvWM3T8OaqA1fWGtT3uQeShC8R/dx58
hWW7+pfxlzFQdOGiMHI2q/l/O/oyP2lSI59OyhjXpfnQYge7vOJX9/oCEkkFRJ9VOQchUeqX2LQQ
YkTjL6+K+gBzu2uFVUN5o3yJh5qTjoQX+b6csaBuVfpBmqXfXAdJ6H8z0ciV7OhDXT3XI03j1SPA
XawVlzHln7sZ3nYbjYLoSb/ZNvcNoRdtgOVQyMkRfEiHQn3Pw0IQYQR73U3dSdz2uW7MlSjAdLmA
Gcst69yZ54cz9m8F+wLUXH+klwEzuhNPYQMQT5/mr+fsuNe5w6rZqiVOyEhnK/kVpkRF0xiSWKD1
F8OvyK37ErJ9zONq6uizfhHjFH8Ku5rBe7rG4GFNNdjA58hUcQP405gKzDxXwYlH9KJ09k561WXr
vTICv5ZhUxFxBQVDt0Ir5j3gI4fW5ih5nsGv21lN1FgWFTc7mYo4w0LbHBa5cHazPKQh/j2jANfi
vFHgW0sT96yUknFghBeKJKGKDR3kfnKd2Cx6MYpqjs/97S7DfiDytNHW8SCBaqxVGXN6bPP2XTTE
nAd6FNk9920+6h6XcWddCipDGCDoR+ERC54ZHg6s2+Lj99vGC9oI6YjWekbkcUOuG9E2NG8yhjhW
n/kSwXImeawnm3wLYZ2XzAsSgDzJRJMIM4savjRBvVyVdht+tW4WkXEjejSIZzQQEfuT69ceCRua
qljejk6sV/hkF3WYtlgpB2s7raTIyzkJwi1G07Bvw3TIvR7utozVgGiKGXlB6k0QnAqBDtR4pXJm
ReL0KAr0WAodMnndZ6AZ4wz9gdTdfTDPd4CJysbyZj0I4uNlrD+clAWV0oPBShNqMy6gMvQRvNo3
gpX2Q0fpaECrBHtF9RwJ+Wpx+eUbljPn3H6KBj6cYsp8tmV16mJaOajW2ugJlJQJBwePRzr6p350
0n1NxbNJx5tKaeHzswgNFy9mviBK1R/qvxH1bR2ZiT5rj3eeFnfm7RsDQVQJpmH5xxWrcQUUGAhp
h7baSTD3O5ugdohb1VdazvXwNBjK4ZMiz/IyeBqIxe5fyHwKYXFeyWUWmnA75qCXd8RVwb2U/WCf
fwAxXUMXTF8jR2lI18lw4pm8I9uNAFBeUo4OT78Sq4NsIUrWRcIvY6YbDw60K9vCTWAURZtVZhDk
Iycd3SLlSbiNdwesCujEhAINthHtC0ENnqzVrmgoYTmIUXXqoH+Myqx99+7cpfUXDls7mSxJd/y3
k9xpU5aY9hleoczZZf48AcJoWK4W1ZWA1wknrhyfZHdiOx9BOM1kqcs7t85Tlf4BDGhpLZ7GHP9l
HM38p3ek60Vv/a1TpSo88SdhWkNy3Bl88j4COy7PN65W2N09nQtzHvGhQp8usBbFBBIfSouoYHQQ
PGnK2J3BeqH76w5zzRx7DhXVT3q/O2SG28fP9D/BeVofqji+AXFnpd5Sk1EdK5q9b/JuaNFFlhlw
nWuJVbnUFv94l2qxoCZknQeaXuCfaxP7ye8w9x1WPot258EywdhLVTOrAP0Z0RdnAEQB0bIdskv4
oLB7uiVz6CX1rJJDpCQFnruDPQnsfewZAyUAHKFlWdiUFd+uFS+zPSunBzzVZ/uKIJHgPD3rchbf
ArFbvnkHJRp1hEy0vbZMDIrBwQkyaLi6ASNGY3uOn0LPVNlqdmuQx13xR81n4PjziRCh4FMLFy+0
6UgJqx0YsBJ//707jUTAGM+FQOUVlyUiicEP50ALFrG7/S0sa1M3apVColnwaxkmSqGv22r1a+hc
R4kTKA+t8VRlfhKjzfmDa/CV1nw2VtjNPXQqN4GANj/BCsNumNTnKN+IZL29iP8+r8K4IgM3J/Bw
4mZO4/zpXo0dtAuAgkNEDvDc2t37cDxuFRg1/8mbcZQkQgWTr8qF+XCpKOosuZZzPJ2CJpVuFFwI
mHLLr7HTNjrB8GlMrbdEhFV7Zh1Sdiv+MAShIMbpsq4+Aqdw0BQv3t5iBkHmMD3JiFTiWeT+jUE3
yAYh/wyTc1W1k3c9zxMFoxhkowykmHPWMXsMYztujhGwJoYDqembhWrsjYQltUSsL0ASVeO/MRdE
ui1ySPTWsK1WGPMtXk7IUwC0IHVMtSmHS/YsIkWW2Kc0knFgmXp6H7P7HhQ2oUc5OFwTVrXREeSG
m68U+UitX7MyMW1gPguRjYfvtwDWYb+rXgSWPseM6rp1UVJkMl+oGA//gNRYJ3GVlZG92R7a/JXV
1THOH2dbdTdOAG3KmvuYDn9HyFLTj0R0bbLNczlijV5IXwbkUescrhzTKj2JCumS232fjsiRybr5
2lnacbPUnSagb4kZYbPnA1Swp8dCer7+3c8nEQ3ptxniR53s24koLlk9cK26qSI7Je7VxkRvtaEj
CyC9XcB5RB1kHAwpOKC9NUMaEnf9NBfJIYHSTUwIRRoynN7wOJRoTZw8ipsInohmnTZyq1elZ69a
SwQbQKRZa4hF5dIYuWiLWhgvi5tHOir/CB8heWRi3ap8mG83qlSaCQRc2ilyWAkJhQWHT1/fr1qD
E9ch8HKASsqCBiv9stLQ6IcVPpnfPnVJxQ8kC2BRtLpbaNYeBZnc6ajgYQj9qiNDNJ+NJ9Jbs5Hp
lDAWH0JRLCm1KE4cLE8IWFUNoPH89KLaE+ziQcLQWhwUp9NFIiYveAsWdgbmtSbWHOIzFOUl5/bb
vKgFlulyhdEBp+pYxwxT5CEqwzJHif/FEVJ3Jd8fC+FDlKPekR1IBJ9HJcGTxiXpscoySQsM765V
vN6LeipWcpcvy/B/FN/HaTXjsK9h4sAY7HUISASDWJW6+W7RBhMgB0PyBWBhN3DEARBDhAjMT7o8
XsdnlvHtwhmkzFDY2puVUvE7da7rhVyheAvUN8v9DJME6WjEgM83lTqrMKIOG9TElE89TzuRzB7q
yZLP9rfLoftsmfh3oaqOcHb9Jfh/s97zX1ndbe8fF/DzUkNbCZbmqBkKw9hBqJAXWL9OuXy9BINx
g4OnYPW+ARjTw4juTl8wcps2jNFUFk/JEW+5z1Jey+2K21tnIm6sc4XPpP7vLhSuD1vLRTxuBCMK
uOFqTI+3ze/w4CeQCGUeLod8EZglev+jK2dnRtWLc0iugTed/6myWrVdrTMrGu84zGwo8e8RrP/5
hnKSrHCbuB1Nm2+TbGxHqQnx7/3RtZ5goLAKlXtlQNOTpB0KFReXKN4JkLal49c9x9YKAo6rqxSj
PtWL9qHWYgnwsc7ljBc9KHK/ZHOeK/tTigyAwiTH4klMLZmX30B6YOUYnwi6vF2tZYiQyskopcTa
pHQKcA2yjDrdeaQUTN19RJd4R31n+5hVUszrF631Un/AZVzIpZKby40ofpgV4XGwq5zG/FW3LJen
dpHQbMb6VzuDAL4vS2QS9WnmKg1Iu9cUQJbC2+idMSlaA/wId9ycohufL09Uev9PRm1GNiYLnqb/
DHprYdngIyzt8+0N3zpbQztOlgAQpEx/cpWjTFJO61bJx+NEWda0qP3mzaYMXaKtpMXCgNg1WvwY
yJs3YxnSkln1+2P1rnCiE6rNBiN2Fw7tV+JWocoQckM5v0G356YfJ05AhsCJZ7eNW+9cgOGNyIQk
N9NU2A10hkw1JfSjLW7hQz1sN0epIw7Lp+Nniw/FJd3sdUCPv3azI7dUF2E8QK9QBQ9+qyMvDGBy
K1lMV+sdV+i1L5Sj6b7JubKmTJ5fbhCsHTEzXZKW3hzugbpzKEYrileWaNc8scA7NYWEpzeo8GHV
I2/YB5e2Ospc0+WQ6mBVunTJNWJWt3eD/9VE7kz7dHMsILdXAHZxCldaCkMzO+iec8pZQqQN4d5q
BWgzaITv+Zy+AbGigkqttipfWvxBhO2CulI+Wc7tjCiE6LcDGeAxthxqRTA94o+Xk10A4o09v6xv
qR0l/vdqnxqK4hX8qWmNxdDjHRs9GP0aDyhEGe/SgvZqa0scvvqNi4z04tuTbwUQPwkKQ8LSzmAP
FDd8Jd9qHfiN0Ry6mra5/zTq46US9jy7pJsi7G9mD5wAtavWmvepP2HM5ZzlMTDAP9T1500fqHcG
rKWE+CmJnhm6F4U3vEGj+qj0phlw0m7GEFDXE74a8YUCcMkwHPfu4Zzdz3dzlHLyEJgeHf3aDBsv
T3Qg+LVC3V8awviMPclYnRu4PPPvI3/UreCbMQiEV+bNieGVDJSCcTqpMu2RRmeRbxZo3c/JEjla
76guY/xSfCHcY5A79eU1TMbIouOrIt+AO36Aeragkje6eG4krD+07sm5ANyJF3ffTiPpdEuprCOo
is3Ewt0Mpof1e/1RfhTBfh6Lp1e1cNQG+pssgVE+ndySLxPLSpGxEr8cu+lDaDM5bcxWiL/AijoB
yY5tV9S+dmVnfWcKYOemBdSqB/2jhPRkWbCRxckDmUhXyzsUjxN367/fobU8iTLOO9euud7vE/I/
IOdJDMm+QjRivVDI2RWvIy7K6ln4vlCryQa1t4zudCiFVIc2raGx6NU3mBjcahio6u8NEUpbprF4
8YdBlOVIRuErWAC2GCS+4Xy39gaP6b8ghWxHdJacGegMSWkkTxVGqyzp7Kfni0xYmaBp9/zDNXLY
oS9mQ59LNphUNstMO8mYVjQNra7ddhn10y59V1Hlsf5Yfq3Hd+a+Rm7gG0yteTLCk06XDOYy96k3
EI0XjqUO04KgOouxBIgZVKOW+CCBlsVV3aEq1sX5cdSUc0oxbDabAvzL38qL2h/G3C1c0YYNW1A/
X7QDhUbOIP1xg+y6iWGybqbHzwXx3f5r5T8s5CbDmozR2DgEn6bg8joNgRcxy5pmbbu266HftJrH
KB4Djy/RkfOrKxIRuyLR+qyDT70kEnl2eAIeHjlyK/LyTYoTVF51sSzoTQzuCWDPx1xpZs9roj4S
sfXrrwrEDrzZj3/Dw/wNbk71PbFU/ieMi93pPiRQVTFmxEkGmRlcPFVvt//g8GUEnSIqzB4qA5FF
9/uoOMRp+gnn5tXnaXaINylmef/6uI+L0hl+OEAE8AnhsAex/jNkRkvyYpjdR0pixxtOo5X0SuJj
uSkAVn1F46suQLhFa8UnVOPQlknLlfET1LGXFMoM15xczy64LafIPLRWqefpjfIKvUnoQwzBnivK
MOTV7g1nqqi78YiCmtpMCrnSvb2R5wIZgOgr2mIsYEtuP+slnyt2hNCXANQRo7AYRwAb29ZhnJz+
AZJMtuIBXuqwMd5RtqxjCUba2al0Ibe2e8brVPc3EA19EmRLfpaomb+B0vEc5A+ZoUUL6JYGNAuH
Ef+RxBxX/nHgG8N+cxhMBqw+efo2v0g0YV6vZw652556aUQyOS2Sm7K4qiCeaK1TIykF1sKIick8
9zZQVpSVaRzgxatIPH9J+IApUErIwUzRD14pjsKMFsAgyQDkA7U90zuEGb2ra/A27I9teff/3Zrb
lXNbRSK+khswCYBtBL5ec67U1Q41qYjyG+LW7U1vUzj6lJr/LBQEWYhclbbfbVg3alnNPnKuETdA
+G1YDjm/kJ+Yk3CZEubV8Dw1OszvnnIUcfCLkaX9aY/PdpMwZKuOgMzDxx5JMkDhPMDDaeRwf9YT
cVOaOxzCToDWCjSTsF/mcXYG/y+esIzd1rqm5giclSpDLQ8wi/fFMnukG+2M4Yomp2P2r4MFTVmA
Du5NuDF0Ta3Bc+FbaK7weFcUp4/vXgmgtUUAr1yxqFOOqYIt6V6zcTvjecxSrUpnm9pz/8AUm6Do
Uss2Scrmt6GNwiZ3ofvvTT1zaBXs5iB4Mq/dZaxNe9HWEmfzVpyITRbGhKryUOPgwIqfO5Wt4XkV
hZprN/6CC98hYp2WykAf8YuTDcP+tIHuJJJ+lDdvbMcOWXXog9Cz8ASfMfXu6j9YtxwwvJ40ZqRu
ubgDqZhhcAWItyr2ZQir9L9aQxa7Ypx+BEbfGzQa6hH5Y8iHjdpoReK71/qCQfW/vz1EE10LIlcI
j24DjQnS6VmXdBU8k2KRegTpdT1pXyvvViIUXdmiTzdC54TvvUVC5L4adDtZTFyFlPYmv8nQeKhO
BgP1c5lbrNhecLBZxDBcyzk/bO+kRJVukLTzsxo83s/aUD/wY5UHF5iZddcdVrPLg2zmKIbk6X/O
a8HHeCpeuLt2+K2f3xN8v3pNdPjXPJ6Y5axyvoP2YDq1GCVGGzrnYh+OVABLPvX3YUJh6/Vgh7JW
BGNWxzHK6NvEZWdpa7XZaa/LswAHrnMYITOczdJRWL0FJintg56LyhH6clJVNVX8OI1s7wzRRmMv
SuXmbYLHuoptpSbjZxpgXcaQ+hbYuULcYKTnsn7yLVVFaN5GODA4qPVp5TsiG0rr47MFS+nH90H7
tFURWTkpZER4SxNbDEP9mriLNKWfFKt/W1RGSZ7Ezzkc/vPxkI/kDt9mx+44JxBrUfAiWc32Ws2h
79R61pc9s5lmBIl0q8Mf45peQgehGRac58G8QTLENa00SKcSa8y7B+YxONVtZfvaELh/LJxtwfGw
W4UllEZ8sjlgJ5JIJzI7W5Dold1/21AEJoSnb2i6SXMrgbk3ta7mFtt9rlE6kRoO7tq2/eU+pr/9
XZm1OAyntrX5xwwA6OX01MhBPnmVSxQ1i27vTtZ9bIj7xDZgEr1wgr85OmxsOJxgJnOZfOJ3H10I
ZlgFffEfg5/YHRFMBSUDP8T8SNHNo9+3DNTHhuTTaPlUoVftMjuPhHv20HrGxHCal0uUn+w5vI6E
DjfRGsqV1gNW3tQI1gtOgT65Yg2bWPUcI1/ZHx1A6p0jK5k94ypQok5e/Ha8M53/3E4M0xLCzKVb
K9F7O8cTKFDXTiFVJ7iTRWrL814Ngeo0UABkOlXt/VMnm1lZu6Q4nTs60Ijp0GZYSIwHS7VcypvS
EERmbFWiKww1O1R58hLQklAABcr/GtxX7W5/GPOaB9Livw8d/KSuheoy/p5+cvNk0a6JMzQ/PS0d
31T7SSJXbjJ9rXyhKNFcMBbuj4b0Tal2TJvSniy3VzZgGbLCXDZ2VBDrl2w5Y0xYlZWQ7rWmYpUT
Wx8DrDzwOZGES1dRD4/BOJRfx3wghpvuwvqeDXs4OtmXVNeQXYHrqjIlguaC0B9ZW3qF5fVkAxOv
3o+zWAEjyIQ+IILhmi9NqLbA1Ix42YTLSPaUCWFjx48LmhIpUk8QbBGGXxk1KGi5Dye2MvChPAD3
KFZbRIlXAAKAuUjQ5acsNvoSbzD341vwAxscGg4Yqt6m/lTv0A4yIu003cYfiL+T7RGMpThtQsNl
7J09MrtLe0qIXad+2JUXmoVrUW+XH3R1K5n1OjIz+gO+miHHZ6Z+BnyTqhI31ukt0Da22mXvmt0X
+IPHrkb8VpSKIIqKcSTXsPCZyUTHg/NJ40IfnkDN1bu2k9KZZaMl/pQMycyzKvXLYpDQANoAYxae
uHJANZGGXDYirFh4Oa7YA/DcjB59mFg66HNwBGD4Ii9nPormayS523//jAgL1lHdFcQoWEHB2GxY
m64WusoY1oTaTX3VYRn1wQbcW8YZyxb5RZC09fKy0s8fuayPrXiNQysCe33JsBWO8vixcEYBYBYu
cxEq5yZNNeN5wrPIh/1GYFr8wruyBfoBFdV+XKIT58UCK2Iajg57or9y5oaQUK2q2JndsTkUo8vp
bG02H3pzZ01uyli2rO7Eu83wokvPk7cnSb6vwiRr2enODCNE2plctvQo9JRpKCpamAsKEk9Y/gZx
mgS7otGj/f3sdG0KA/Vr14qrlq70c6tYrf23N0vapFKHJ/M7D6A9Fv9hZBFLST4DSeSdsFE8/4+K
DbMMoli+9mrS/jwl+Zye/7KAS2wjeQEBK6UlFWdEQmsbZDfhT0n1Hi1EKbDJGZXpOVliRY0JDo+v
cqvrew1eFAHvA5SazqRRpmue9aVdqr6hHuhXiNan9hok4CwBsrfYhDvDtcSl1D2eCDJyxtatv6xz
13ZY7Y0tw+45t/MukXzgp8JlDrm8V3duegWbK8w7f1YS2ML9Msws41C8qmy4e0N8Myt+BAkQs4kI
yIQLMp4FiGdimWlLWrVDwMmrvBhEUuGX19YNYdz29OvQgcUGz9C29vTAPj15SfRmCgEqKOojo7cF
MgIEJM1DaOa0hMAvSS7hTUh8MJPzbrcy64YQpJf3B+cZFaM6DpHog0YdrTnU8uDx7D7sR2Ua2bYf
VBlEsbYDiMZOyxbhasBQ+0ccpKEf2BudPXmNIUuZEfDR03bub6UU+HNdJ/aqwbgIgh3fBwzJBgSt
kNdxNzwUwsKK9qwcL26B/QXQsftYlv3ZhmTYEu474MxIgXTyDIDsyZpq+QCRDogIjBK4hgBGbgsR
LNZfBFgKDYNoSQSB7p0k838LizWclo1ZMURKzK2D+O5/E5BwkbHODG2Zfe4XViUz3GSfAK8dEBHK
9tdJ+RqlGo+o56aW5uoCjUogmfjsbeDRFPt4KW/4cNlT4dipey0F4h/p+MOUMSeozJFad+3L3zZk
96pDbA+e7gSvMF0P3HEn40co88QjPDKdkLdueHjrm0jVw9YAYw3/3LSA0Y2B6HujHiRC4Wp5+ejn
W6IBwqY26M1pFIXLaDlEA5QIc4SM5Ej8plnTFLVZvBMukw9zF+vh3NP74hT8AM7XpselGlGBxfdx
YOIvukMbks52qvfJKTdptBMP3YKCAdRIl84zkfwvdXm1OdVKePUaHkKkMWwxJT/qtJ6qwvMUmqnA
cBWt/B1fka7TsQ5Oh9JPk2YMNWAw5hNdiQFJ6hGLsE3ENLIszW67SZJLzB5D1rE/L3kp1kCxVbWV
wibjo/NfQQ0PBhmuSDm5XSCcGFbIkZv4DQLSdESTZjgnF33xxaY8hpk42jdIHq03LlqF/xJ7XR1u
/akU1JyiDBVPhAj8AUIdZurYyZ4H+8jM1OOkH9aiXRU9oQLI4+6n3+67y2fOgfm2ylY3MnK5Zuca
AlwKWabVcY8oZ3VzsScMpcyy9abJV+zZ3Zif1gbL+zwRMg4r5wpB3vUDhsOFTyurj2WQb1u4zhmO
hDj+Jzjq7xF6E+xfZhOHMOrebFjR5den+Ma8SaZcMZeFkhvNcj/qeuaXbeed4huI77by0B7Wu5nD
PylUOQlKkTG8nngN/SJBW+r61B9kUfhovQpge9Uz0Ux3GXKjyPxcV8OmR7WGHyRJbHqlPsSmOFAs
ekdEINyPlYjTN4ZXQ1wDYN0gFaTr3bhcM0xr0I8ewrBQcc0ZfRg19eBdDCYEloOhi8Gop7abIafv
1E2MBt1Q94Q9r0s3naLqSRCom9OlyWR9rRNtsQ6ZTysYc/wqJf3SHVtzWQmqDfWGa3zkp7lUlkg9
Dvn/3VarbObZSE6JUqRI+FZkrs/p6Q9P/s7jXgiJS4Gq/q0t/ZWiHyfZqjZjwYIXSRVk76xNOyP8
SOAeVVK9EHx5B/rMBBASjDaWxWyU/AMzjgLelvUky8cfq1ZKG4NykZvTrwQAwbWYPcRORmh7GfpO
zP5f2Lh+uQwBd8MPJf8edDKmmzhqUsdJg/8eAHw83p9GaoZLEW+ge1a8+yWLblhhk/7t+CNcNI3d
UYf1e13E5q6BlWr42gx0ljse1+/YaiGE2x1ZWrCXcf8K27VaTZBRkkNWKNFGJBFA1k0xDFMD2f4I
xFgPcCKQrFj2qh97gibfNVSKpx97dg93NRma4l0BTruye9+WsMp0sjBzf2xegPJ0tUqs3LfZpAwf
WntcFLe2/pZwobXNyE6zMAZy9sEeA/lmSsJBbk8ex7c2PN37VFotPGVRdbKn0EyEKvVmragcJW/3
kN7ZmKd8pEyq+gT9MoX4k9EU1+p76EtC4B4/yM3IHyI1yViQrcKfgkIXQ2zfU0e4bzmzUssu2CMI
pVTFGcT7idbu1gekqWBQ0dpGPFB7dq2tQ7Ri090WRCrVXruYeElSEStDOMFba+HFwWYXvU095POO
/KM+1TexgvkyTEKd803Z2uYI0NKTh+lTv9hdAx2wUy5ExeFPScD/tEVyTkmdoHiAOAKtPVm6aVI2
KnIXJGTQY88IaGinhTxEMt3RYOlNSHdFON4szNSH/GnE+Qdp+Rd/kNaioansekIhUOpNbWvpzwCv
QJhwoF48FYKDWb81rR52p/nuho18i0T0ieahJjntoNk9RCX3vKTcUdwdKhuHyRYwB0iTCDeyeurV
YC7l9f4TeWwg8zmLYHkASQOn3NX70uq3RvsSvo53S+6dgp4WmQZpBZV2sO/gpRKnOJfe5pGbBY8x
LevrTXr3jbIOqm4tNlobDq0c0AEXcrzzzO4BvUF7fS9hSVT6ih3G6qv6feFobPQKvQ9ckKKmNwQH
KUSNT91a0q3divxN9yq8YexUm4ltcnbQNpZBKxEYBK5faAgDrSykKpYu118sAMa92Qrt5lq6Xbzx
GXhD8+uUU9F0bfNlWzmAy3MSZdASUDUeve/oi8LQ3hRCmpT+8pa4PUNFoJNh4FuZjm5N8v57d4VR
E48fClGX1yO0nDBE9HtFe+F0pcUPELnjwzahRQWsQuS4w4E9KfEIhyClAR+sNS8e/kyUHPSAvRcs
5hHGu9VmSPL/4D0i1NTjQxnSmTVrwH7ruqKP+REDIl7sT0FX+zTxiHPWrxPp68TOxSZEXXwnl9j6
g80YtQQET0ode+tZeyZUSrp6UMxa97/2DILaH7O/AzAQn5He2c2Y1lnTjfifZsl8jiWCYexgRY12
dG5nrPCaEjvWZQZljqdMbnzUmpQ8kMP1doggsDIwV+hcHbcNh4FlYBPfobaa3xzIIOCKqtWKHrju
JiiDoDjlmVnJc8QRzW+PowhIIEwdcow8le8Mr/t4xo5TGhS+omDf3c8D40NTCA4d48XPjOGqzuwD
GqXacRh8JKHpmreUwq0/f6J6TMAcwO4I8z1HEz39gVkfheitZwECoRyckDusi/WCBZTeEsoc6vqO
I7LBD2HTEO6K6bL/pvUaX3b6B/ZIfTBEIbswoQh6HEhFWPRuWgMlndqriBY7kgjfrA93TYrHY7Uo
iYpbpEE7lEnEBiDgwKy9c27jYB5qRCRMfw8J9v6l1n+EP0g2+089OPcGgXFW4efjo8K7MoYPPybI
fdw0Q1YK3C7hH9CxZra9r3uzLFyyY1vHy3VDBdPOOSPrvfVQB4gEZ1SC0NSf80oneIrOMRTy+b7y
ZfJ+SwZTNhzPyuUzaYvKjeRMB27uhiJ8ls/bXgzr1+UW88D9Yyubli+m8CiVHLA5yJH3Rp9UJYdI
rbC+kReG5+g4RqFL+fP4K7GImfpm/KoW8Su6xyYkt88NRi+ByXOjpf7HqX2JSK3cMOdqERoCoyaw
vO2jzxR7dLapyBYizRy8SdgHH138vckc51ahvafgjCDTuK3xm7XwA6Vo/8y2B6MoHcK3cAHrSURa
aLUb+2IiGqcaFGa6KKgbAq59tu2hh2kePLOA3uHNcGul2vd2upe42gCcMt81dUnwpTIZze59ETUN
VsLHKEIyjUVy9pSPm8K16GNZ7Kw7nclhMJs5xMWPoYVgyaJQ4iAjA1usZDbjKvSNgNejs29YVlfv
VjvixmxGSJG+gmqVxa2xaYlSWee7w0uAJTyCoiOeytLoGkFH11uEyQNNaigLVltKjnRLKIE32Sbi
jOWdgFQU0ZZ3iDdTJoWDW18C7dfvZ+4316Tisz7/fbatRlWeq0IBKQWAxIidIJTCsLWoo8PoiCu/
tXtYEsmn05kxL89gB4qdv4Zpvl0sGByiAtbcez3ohWKkvfZlW5IRjNUYfGaCV5OF4IsXoSCo7qbY
HTaM5IdPGMDzD892/SV4pcXHykv5SLVDap/WjkbkP/YCl0qRSe9xFZ+VMJiXo+QRHuFjH+cVwM7/
/SPCoLSc2SQmScXr6yvkq/ZkvtQRFs422KkmeUJQGMKzW1F8iKijl+3QIx0/knkBjm11hL50YLfX
opMlccDinT5gRih4Qm+GluxwcGxMKepHIuEjSjLNTgFOYjQ/tDSssaEYTYuQZfi4TxkH9ZYjpxCl
rQpoNW2AfUPky0u2K+CPbGaYKnvgE0OUNl0A9nE0e49R1Wn2vZ/a3iM/J2jNyjPlFaU7xHZ2iIzm
Iln1KfASUBGUDpYwnxdj6bz2NXOo8kXNrXwDHt2DLg75aOdz+k5zClFWCofukjLgTigTV6NxeeJk
8WW0aivle6615rPG5k69lxo5AbDR/UeZp0pwnys71oRUK9pHe0GduN8awwRN765fJQ6oALVjMhzy
CHTubE6MaNjJKl3ZUGGQXsfTGr0dpHyqaBgm0zEd0PNTnxIlvkvw4m2oj6arlK1uQJ4vY1ettCvx
GYMJl/JFOiB/4zt36EYJ+kFcrry4MCe8Z8IIO5Zhj+tyi/t+5GGMPDU+ctMoSFUaFV2jlssdU0Cv
XNpCiLhWzVdbxivpQ7//CSPSEaHgg6njHE+2rrwW984Jf+qQ2eO21xcfmt7PNy046zBPGi9wHD0p
l98WqeCng+fbxDr2tGDH7JvMPHbpG8C6b7F2la8lIYU1bVJeGEtY8vWGi2KHP78EcpxdTs4iHc2a
hGRDgYXcAB9S+iSKicvDla7LtLVuce4EXudLtIsRSoXxfkDvLiq4ve0YgFp7/3aOlz3afTpEssaG
xN/lvB3T6UwIzTyfdhy5SK6Y7AylAoP6ZJP/vjE+gd29OgeVgpLWnLrJ09zw4PyL2BTSYGNmy0hO
yfXe8BCR5gjFrsZrCmzf+2YLVS+8ywdHyFgXoKOOgO04SNmsE2FGqgxAmppquYxjMgLBtT/LXzcm
AZG27ewJRRWYi5jTNVFDOrN8G46sYezRMoyN+mX+RnDp4z06Q3k0uPV3F2poIS+UEFcawZ9Sxrda
pYEWGG+mnS3ocxnl6/KuN8XgprSZL9jFSf5lXwDmQSkjsdQQn9r5PALBMKFIOqdC28R9dCuuNIwW
+cYXJlC7OpDbk7aOSCoSKWr1BvrWj2n/XDBhCDus+xU/QfLYfkFupjliOUCnPowrc0Z+Mn72jPsa
3uvCEroNFF1H6VMPEI/66q8FVhY74azsMmn/yRTs+T7liszBlDirx5rqAyU2TPaZ5+YFKoGXFCul
atOpbBBdlravnnpiR+qBR+oYipDLp8QThfBs2Rv//e580DA0wCAHmMu220TULWhSrnkj38GnJRH2
XUSjrui9CCzYbxjeMd1bYrP5NLQYgHIPFx7eFfmv4ENn3BUXWN/wxeRCpc1arcQYBNH04S+j4vr0
Dw2yPOF8igK6ze+KHrqX2SaHs+1nR/T3wzpf0x3Oz7ZQnIEEyrY0Ves9P2EJPRGH/79wtsXEDT8G
HHSU9WLk88AESeR+Nlk9fC8Ka8FZar0YF7uxL03VBJkcIkaUFoRY2ua0W6GvnwXE6V98EvCAuGof
argMpJ1OP2EfahYr2e03wofyE0fqGFRFcZ59PKjl/9H34MIFHmjdjvgDczDUeAZRnSjy1Kw5c34X
fYcy+6T/Q2Aca6+qAaaWo5N1MkDrgj+otMix5mXL3/FCMrGwElg+h5e2wqQmEjvbA7YAr1tiIGWu
Uj2KAl6c35vZEPpbam+tF6wpxAV+0cfpJUuen5nsHxUiXDjUSBtPxSpwWd7bcYADPx904DmBa1Ym
1euwMFiypjqzZx5cfIfys/wLNWqUvPT8aWeJtQYctB9FfgmYfJtw7SUbbXyL4d5Iw1mec6GImnOg
tKc1aCLwJlyA37TRa6wolMvuX2ADAoJpxcfSwqewgNp61CC0T790HkVmtbf853OIK4yQjpT0kT6Y
3T0K1noG2lFlu4MmDZCzatW6vy7c8LYDUef9YnWB+X0PRj1s/8W9T5go2nrJsHUMfqExKLc6DWfp
wK6va7EKS5js5XyIxMMp1LSORtbex37HztTf9IEjqWzyOQIPABNvNe7H4TfDJLIsus1pkGDW3YCy
vxBIVvnYr/tkMxiQtHVc7u2MvKvG0qfgwkCGgr3ureWmWbej5rnryaqvNDx/zB4nkTTD4No/iaOv
uCdbkLFg9HYD2UQgWfDkWjJYLTqCZXwcxVUzXbG1e34urdbSknZ9hnvnhxRn/VhAl0q3yXoN9EBB
tcn2J15O9Jzh6c3YuPUlKfXwMucBh4Q/1Ntc0a/B0P+u3Ni4rZiRwqlUxWENR/YbX0mquwiME27y
lkbUtxrmGUposnx9zIs2JjJI/ehSUtA295efxw3w2wicPlOgLTvn5OUEO/MzD3T6edLSKU3LTT1N
wrqyI1q5o69ZS05gmzD8fN60236T/iMD2PijBeKGMokcmrgFEq8ZylOoGq3994AVFw+Nx2NZcViw
CnmV/iXYls+bXNqZ+iQLz5GTUHrkxBSxsAuQvsV6Vo1RcIrh6mdah4S89Pa12djwq018mZcxYvcU
c1K1b1y7k6r54VPFES9B8sAeZDyZGqOCngBXL56R9ZF0wQqwRECREhdR3zEdO0Nold1x+1+W4utE
aoMcpaeahgX6OVjKbUz8Ob4u5XwD1rz5El8+aGCwOz/159KtLxQonW2FohuEni16yn8UpKKud98Y
d7+dnG83O05+l91Se0Sofxf1p7/kGqcWIhkjmNvA4qeAH3R35srbWMJpEvBhkhZraAXj/I2a/ldw
RBAIgDiqiE8Ladz3EdSqBiLCBMCDNUpFjqUgEP1qATIe/vdYNiT2pj2ZAVL+sfa9+AQ/sW5APe+N
0cuTN+Mp7rY52N2l3K1VPxCTnpQGPItx5q0GSYuTfOVKx9LJAYPy5aYCCG6YX32fsh2lV9ZExVA1
MS23skE0hvCDulLg3TCTTBBo/nLMqxucDwDHPig4yVyXRgu7nR/g5zgiN5LS06Bubj3PIy+CbF5E
7PqWzLxTSR0jSnTW6BPViHmyrBaJxdgfeI8i4f4hBqnnbAkVOJs42oZcANmGWm/+VLfPsMsxVeM2
9VsGRZOSwMkRECIBBKr9tCpA3XTKSAfxkn9QMfRwz1x/w1F0C3e2ugwsT01L+xgh6wrikDTjsVLB
yEla+luFvcZJX49CwglARADm5ORMwogR6osZ3kBxXcWG6dbq3u1AVJCX9zLccHPZGNH4OdMNkcoR
Lc31EDb9DApUEEPS3D7Ze5gSKTNc2zUrSoTlj42iJK3wU6KmCDqJfeKfJG6kZSCgdt4kcM6poEiF
FhlDsIE9Ghz+65Hnd0B2tAIbOyY+iXHEiqERnvqqtwjaXP9dOxnLXioojCSV5V7pbU3GC8wk+X/x
z4xj8QLLy3tlbUqYKd0XlzpviFlc4cAeMiQwg5AIVOhzn8gOOZ9msgP6ryDza+5ocyHa+5PDvdPH
6AaZcTI5ISuvpcq8AfOTAk9cz6eoFZZM5FuoUvyQd/iJ8mgkvitC5TkDUulu8qI18ZcUz4UKSSBF
SHda2AqskhoqosgHbTL3Wev1fVIfoHSpH03FFbfnIY7AnDqAGf8DiKJbaTJXWJPUyhcQD+6/02zA
nRov0USFbpQu7GXxXqTYAimQDOVl+CQTqE9jynOcD5Y1uxZo/e+8c1CYfOhkRjQxFT2hZCmPJM5e
KAXpuCSfNLkLyMtlA1jUDq3bjmhDVrOWaZEH9eAK9RsX1noR/wHxkb1ebzIrut2WUiOdED4OF4rI
/mLs3GcztEmH8m7pVyhCwdfQ5QeDfU4Pp6fve2xUfgQqI6rduhkiilyLVfuvS46SPSKmyZm8Yi+R
CaNShUNEOLH2WYGkwxv3i/ZaoBiaPfkaCFjO1bY/ZdZiDoy2f6vdV2yENctbDr+XNsxZ+lHex1kZ
+oL0XOc0gK08fzdyztLE/nFTZsek41Jgg9Alc71oV6Z8s9Zvde3/akrgqqEBoqxf7wRPMTOnEuPp
iNxdeB4KNVv5q9Fev0b2doIJLKOQulw3J9eWy7ee5iwLvVVdhDWMYoPb70dDU9wk9XGzt12q+JnS
5YwJ7EFoO5JKbXNEAfyGCh8agJxZL4Tn1txJqllBq2tL+k+ycdxUnS7riBSMD6ebeTY9YiyWQBMJ
k2EoPvpWIxNQByPOlMQxeDhp2mn5i9++atCGkZfV48BmD3U4BjDcvQPguSW8WOxSj8aKaPyZEByn
7KKDjFFyaiecci8j0Nx1781unkhVG5a8lRFQSGf08x8mL8/2yVw3We6RppmSfk1mgfsiuQ3WIqCv
6tv6c1N3pBtUJZyY9e0TG5c0JEE/LZFzY6AOszQVTvoxfPCnrz11tDzqxCw154bsz2VUEEVL7o2h
q+Cf6tGhfB98Hs5o+fXgirN3YrBVqHSgIjdi3oabKyvswrDcgxtNkqYp9ZXcTB42tiS9uJyo/2PF
fnnqyTlgaBDmorO2htCRGn1uUN+5s+E5ZTEyRyJ9q4TmRsnIGTTPXg2EmKTCedbsEitjAigKEDZV
KtlccgB/1/rvKt9o9HyEyBda/BRLReWXLQtIrrHOHdTNihzg9NmZtfWEg0iK0UFle0JcIJ8y02PJ
4NJDpTIA/ip9wWTCw5w7tn/qJMb5mZmcrua0wUcFHHQf+5qqw8+bzS2s70UsN+PvaqV3RiljF+MQ
iaUmySB6pG63uZ9fbuMeuV1UQhpFoPPcGjwoeD+UuzxTABn0E+uP3jeD24dmN5wo5f/Szxegya7y
7WG8x1Ws3Y4z24EEINb0ZAnRIqAxnlYBfhUQH0T2UAHQiuVwfhe4KqQmkcumUmpg5qXBqiQxeR2u
sZ0OONWLt8EuYR8LG97xvyB/mPUtvWO3us0zWanTK0KECJNaSlsT1CrbL0EEN2QKwP3uHkVxPgfi
PF9K7IDqWuFjzyPIPYerE7RHiYLjypPWFovOJSsAtpF28x7doJ0mWZFylGWzP6gxlJq+mRJZnggE
iWu0qjc4OTVwiA++VrDt3C9ouKkzmKtJ5mMDMsYsfe9/HWHyoexM7kQfHf0aZrzr8gCM/1C4OdJY
lvXkFq6zuYKk47zyDVELCVhU2g93oQNaGfhcX9iOfQQM8y1DqaBVQCDUJVv5a7xBB5xXijniaT2Q
UQQYUnlFcY9G8SKVuE4Z4PWBoYQbIedfygnfIk9EOse8y/V14vdMSzDBBY2k2VgdlhS8YgnGvKlK
EsGPv7Hw5cZaXJkVmbXOu8UH85mULmCd/cT+wHc84q08/Dp0WSeWQZDfrDIHKKZ1yQIp6b/Uyoad
RQ410Aqq5xetNUo5cTa43iIV6RbmKPoTCHrxOkRfF7y0lcsXQVRJoV0IAuc+Yi5yQ8Wn8H0YMWr4
oszGrzk2qeABrJnvYFQ1enewv1R1pPRTVy1E9Mc8BWQO1GANRur1SVDKdiVJTTHhm83uqw1DLezO
UrlFu2U2CbBdHhVzhC5eAdH0cq8Fh9imHNNnW+pmTqt16HK7Xcnx3duHudcYistNXRhdV1lRzgaf
JbMorjxwXJDoUvk46T4lglKHlY+vxOIxb9pmXG9OqsE9JHcYzYOJuqGVE4MM1TsINfsBXnzNRYtV
60uKTZnZ9rp/+2iTguJp2xqNn6oMt/H0qmcq4avxEan2A8CbMPT6Yseaw+ZFv/JpoQ06tsq43NLy
IEjq0EfADEzuVvwrhUPDGiwdqRv5BwKkyarJzzI0r5/JflgKcl9nkBfKSvx9s5d9FIGjYX3GCubk
AuJV2iNnlbi77Yg5fyGNtzhG2+4ORHSChTVgdaTMU0BwmRka3l1/hOtOM3Kc4uJ5O2IeDKmkYdDF
MSxa44E+QjP0OaPBhiIIk0hKhMTKYr2Ee2y+oaU1npJ9IIQRyvzZ/4RSaJ/icUrQLgtL+/ptkBm9
J7c+5CVDxOgZz3yC1JfiEQ14bVUn/5BOdJGRxCvfl3F1n8idNArjKkTGQmdzOHYCOyGZEXY99fUy
eYdpIE8kh7Ep+g+CNHsxy8YepIzxtMDaJqnATE0t+QFSKRN+QiRzColpp5wGMGHIONPhm+o3yP0T
PF/VeRmZ2JteP7WK8Lb3r7NyEEGJVKhEM22mS1uIw3qHbQRKwZNWy/1RKlwaPLa3w2pYTfLO74LL
MNsK7ZX6/4LWCjNtrtLdVgRx15zqYZaN/AA7Jhfxh4PDC18cD8ki2N/wQyYJ2Xp8V8IkLbEev9Pd
bwHCSODwSVhWEKwLcrpTx+kKf5R9B9or0IXMV14lW/CAxXNgo4yfGdtK4ZMmksPo1afwqJVDOh9e
SeRfaoRZRRe53bbLo5+nu/u6BN6Gy2S7pg19rnC3yE0HrnWFS0EU12UOuor55gqxPgGIc1DOvLqS
jLx3DUgFfZETKQqByL0920PoTwDseH5yGlomBujlMRnQf8H0rGFNcT3qqMoGecUENQJkU2f3S4k9
L2lpLbhBrBG8BpNn2TeNcyJf1N6iGUBbaKTel08tMaiJEMgcKZSydpaaUPj4wNeuBcpOMsL/bykW
xqRW5nks9HNa0w5QI9NdkVYp+Yh5P7nWOZDGMcIEN3M5cExdyS1/qATl+E/KxiWFs0qVNoJhIzor
+QCOLd0GY/yNI3jVsA9ZkP96SJp1ifzSLWwXO+1YK6CjvJJ0lsBGbVqsYT+LqLsPVWNXDmBY57Rt
WSJxVEvSU22YR1CitepDoYxks0EAfpQNsO8mZ1eS3TkVW4gaIHSVYzGhd4HdaYslFjP3LhDJcu7A
nO8LngGtyPiH5mlMVYc3osAzOKEJiaqM/f3la/X1uccjXsifM35gcIYyFgJje6ZCCff3eVOl6r3D
NXg0w4DUcERYqeySOQlB2fNlUYuRqUrnUJieUP0wO6QiZvpagY2jBXzHcH5r/38Q0w61sIXMYFa5
x9tom2jCqoHJ8LKoc5XTMOIlVceGF5R7wLv4r99OKbAlhY3lZFpxrJ7BhfLnHSXxxmdOUrJnS+2N
pk/OAgzKyijSxOyn09jgxQgQzvTtBO5TXnIv5c/93/BHZboRuMuxYOuazsgR6lesuQerCkHMwQKk
7Bpi8f8ONsysFnrKtKzDKPYUByyqTXk3NHKZNUHi1phKyDTBPnLnwqR/T9mmccdllacRgjX5hywq
Bwp0wail58Yjo9Slr8NRH0IV590wetGyKnzSDi8qEnz8F9RxxksAoygyu0acNniyrz56Fn80234T
cmcyoHpfyQB/o9nH2L2Mqv2JumekUdSPWqc+22bRHxPJ6VA4XkAKTEQjoqUnxFVGsU+AvyjitLc3
qjbNgTWfUvOBunStugKZ/wdphz0A0sNL4JJkIfm68yKGaCeL1gRVMPTrwzlRXrkZLHGl4I1bEGqY
oR0QbiM20t/8Kr04i/LY0+GqHcY+EOaV21viE4Y8nY0PnVLt5R3X7bHj/+tfSz4NJ1Brp+f9plTC
vHor2OwqCiWLobo6yMUrEzIYuCADoOX38Xt9FG/XDjRAfFz4T/x1INyT9i+5WMjOxlF3OKv1GZ4l
B9Zuirig2R0DayvKphRYTddE7iUjjXoQxddYIbziMsAOGvdwjg7npUpVwKOABATribZkTy8nkl2U
kyk9gF1bLoogyFuhOcpQLsAeB15+UufbNzFG5i0z9HaGDSPZchiKArofbddp/pf4lz34odfv+19q
kQSj+5LfAEpQaSjQ2JbCtd1PRWAkHNaI/j54w7Yq0xiE9DCjSqbB0AXrTzNVgprM9a5c/DsXOXxu
HTXI+ekCeUP8iz5lDE2PDwYhoE3fMxYw+dR6Kwer7s/oYqC0Y885aoSYQwE7jbC/hgpvyPF5CPc6
21xnis+80fiUDvELg/i742pKdEUuQ5zAH7twEEmJ5hKSni5veZeUQn6v16dhuydKaf25Vs01L/bO
jUUs8S1E2V/N+3GILOPCar5TJ+a8GJieCaaHZZBx9pkRnOBb+4u7BC1VrqJu+fB1jY/RiOUhyMBX
i2S/+ca9WABUoPM8uMJ8gnPY1oy6ntBL8uCio0kQWrvE0jJCRue2OOg5PZ2KJzUQtXAnGGpby3wu
IyoZCLEQfZJkm+MxIDVAFCb394Uy06ANe031hafV/PlKBpAnbAo9k29wgZl2i8Bu1QKuWCS0a4LS
2LRcMyqxXzGb+dAvn/Xo21MY8Tv8D9xQkbVXBSk4m91akfrr/z3TRoyv0u/HfqwKWDjl4rQBRSb+
1uHoPucff9sCwdysSZB7ejO/6brUUuFNrgjhpiAviMSlntAenraT5fHGcToWE/VZoQA/kLLkV+bG
Ju/ZvyoBeWadgGQ384lIZT5vRifQAv+KVC1LQwmpOWJ2OYOT/rF9dgJWi0f7qFxiQKe1XUxaNNq7
VqowRjdOuoIbNVhZV/8ms6iJujcDwjE1K9gcDGvPsfmjLB033GwybZ+ec3HWJpdSvxR5QEmp0ZaD
xQ+JEJ5GW66ewlr7gVQCNLLjgWg/DI3Kyw/pF1kPRTY9triw0c2rLr9L7BLajzdzu+j57hV3hf3O
PitlV/ry3BFSKuYFKtabistgoTOB3wygNPhEhooGKzZKn/f8BHHpV97fHg4hreZs/knetZldJQRp
wLpIMtt9SKc05fX3vjwlzgWYeIFpFPlafPHI9E8JBwFWYAYA02O40grV9nyUtNfDHx08l8rdQx9j
+I5Vva8j9Xa2sOxAaxB8G+ivYLapz4BmYxsReP1CEVAM+NdDLNzgxPouJ5p+6Bz1L8FsDolzYRMe
nZFtKq3nnp/fcCmBLHfVLnXInQBlJQEuwdXdOzmdKg2oj2PsR2dPCTiwUG7y62RRYi19+Cnn2e+a
4exefFkTw0hZ80uXgt+Sc83z4coAjlkPeKy3J4yKYT/iC7M0cyLxCV1Ho9UhQObxeEZJy9w6Fp35
L40sOVWn1nSEfZgUpLmvIedaszEtPPqXYzGHIlzBiBeQfJ6EXN1+EOY6vJZjl0RQkvfcKpyRVVY8
/jiPXtagyZ7K/ssPiReplfLbRo7iy/ENUT/MZIgWFC8ZHF913OHY6T8wNXIVPUBbumq/44PDl8Ov
e2qj2b6aFCev8fNYxnFstvKEby7z33DTT7TtBcLNZ7cF9YMZWbuElz8P79ZQ0nNcl76Dg3mE0o9j
LTIJpWvgQl6gDRtpijX0iQFaIPkdXAANZlaCX8WuNG2Y3OT3XHRupt6lyrs9Fq5g9PciAca6xxBB
qdPioPayEq+Mq7RsKwbnyWno3f93umqCH5SDkJEhWxwZurf4cjWNZeVG/cEqRnf5FpDFsSX89/aR
NOwMHjoZV6o7lxrM4KxFL+fHvq5hX59D3dCN0PdQKHODIXvWA+Q5XgqRRVogiiHF0dFWCXYwNs4h
BjyR+rGJBnAbx9Ot6G5Zlmfufv/LlDTzW/5YbBMc+eWGcZVlULOWOP7eAjJfDmQYZoREg8Yw6Vei
Y0PVXVv1BYpMwrVZ/WmKUl1s9RDDbFaEOc/6Gd8krGPbH9uJ8rUGbeVkEQ/qz6LmJ5XDHL0GgObr
3YNjmX5cfw/8zsp2RHUAVycXwroPmXyjg0lAm9qq36+MakntAk+8zqcpYoNKGi9O+G+74d5WgUs7
2tfxs9v75sq05bDIVdH7WU0lmoCWE/5h2cO2KimGGP6KSfzVHZylsMwlwYUL0cI/5EZfvaV9QejH
lG9o9nxkH6xQLOUBewdDhUp4xJwom519RvBT0XjdI6o6oovLyXVx7BGp2ini/pgX+uGDMYhJDDCJ
o8pklFzxKO8EkKvsIu00woNMElzmFksD6J36WCPjWgjiwHfbK58zPQYCdi5Dk+HnqHb/oxPqcf4X
O6WNb1KCHRyUuFA37xTeIpLVg+cPXYyMt5mhklxPCFUbRWMkE+Cxwlc+VGrFBxhFDbwEUHUPs7NU
yteivUcJ5ZMKsCM0hiJ2GLVgVshws02TwS6dOLcdr6Xm08Xk70Q++pasmG3B1K5PlM3dTlwg4lvd
zdvEaiN13aug7pq0Ab4IS0jCtprlq90t0TlJQJLcysw2xHdAJHzmWZHxAhhLTMMZR+/IZYZKPN53
3Qmh9ZFPf45D80QL5j29ALzJhP5cWD+WGdh+jRTtixD1LsMf5qgdBqnlte//C2U7LtgZp/qWYWc/
WWNvNnFGarDdkVcrkYVky7p+oUVx1zmENbWf8rg199S4NSXckZ5420O3KhahmbPUiNAqFNPn60s/
rPQ9ggiIZlAi+AzBWOPeUIKl2hMjqdBCuj38hHY9FLCg6zoDNBlkrIsi1KtkKzBnyqzTKRPtySKV
WK4zFJA7lAj2mDmm2mDJKHVsjTuycI99q4M5nsok9SlXGchYD0aT5B5uZEQEL4uV18xVIi+a4jOt
tALskavdRNixbkDDQ/sqissxQAPANLA0hsINK8XUzuKIDLYxq/xqiSU85copnAhHRSFukKoBI8l8
ykDWR/AUjfALxt5BU8jO6F9OZ02iWgsXCjY99sIb2k8cNqiu80Sj/XxdaqyWy0QSg1xnfgDLrcOF
VFj1vJ4db1paqOA59xd3pttsvJoke+XSnPb3qzPj47p19ODK7pVjDy2/ilGouJ1gXIiGh+mKDD5u
IWEH9Zvfej5QF9qwFjLPeacuJvbvd3Wqv/JKQuJAs1yxbax/7CgTs/ZrEj2319nULJbaaOSikazV
E2wlFIjEM3aAookMeAOozBFCAw+rEwF//H81Lr0bMHDU5sPth9z6pt63Ps3H44nSAIb46ZVAFr0k
Mn800XK3V2UKvV2k9cBuq1f9kh7JEaSGerKXzFD2MEySKD4VZ5aWMOEaa71MkANisPqRbYXSdW3O
aIsP73o47SG3arZ3aaOAaoBPZZQC1CvchsogRiO1nbdiGGcRaewQXbsUhrHnq3q7MG/5tq7J2C6c
afKPO+9Ei7kmTflhKKDRWAlQxeRx3iqqhycA0lqpOTtkKvGXQyu+M5YpQVm5HEgk8SluUQFC099d
cITp+SsvmptHP245Qk2PASlNpgr4Oh/DI8xD1g0V0IlfBPmwAq1gR54Dtflwgjwqt8MDY+ejZMoJ
gw3+OXYJxIi2XV/0tpPSTRSXElLj6RX845lsU9G4/V3AqVF5Fwlgn76pNDH47XKiyUCMbyB3V7S1
I2yFONDIJIjfXAyOMywm/KmadqeetISyJh05UBAzkUMs1GOUNn0grgkJmT4SmBh2eja6x5bMyQC4
s/0WpEex9WUzSGchBMxp3IVVewh35Um6rWhgkwMO+WF+J1sseEJ21kJazHinoziHvTdXcvjuhx2U
OP6UxLrT4XxsQWiXrVILyULeLyr6vRp51n8JbSwt2ft8vQUX6jUzV9byuy60pJauuAEb58AJHEI9
c3SKSrpFv30WW6Oet8yRKB1HBDcbmX5ngi6P0KhH064GldsBAvTI1ZxtbuClP6WKVyRTd6DIyVNx
y/LtRM2Dc6wwTKawOBo5uzyUwmq8Tw7BiXE4uRQDyvz5FR/DTR4NaKb0cajW5CTsVJ1vFjlaDafc
Hej1a7ta9/Pwoo9uLIFszuyenpMJ8WxugYbLMomQjuUjgi0oZ+LtE4jRFakJ5st3Yxh6WGy7uU1u
nKY32B41Jncm6mpAxU9RbPWjk3hgdfevhafqZqYbiHzMJmAmeSbQ+xhX5xQZc+TquUP1RflYm7Sb
cmTvDhqE91gI74KGh6PPtlGfyjQj6vrWjVifXHgIdm2TCF66Z80KMAvLpbIbkkcVaYeete6bkES7
ogPC7FcEMILENL8jzmpDryW2adz5MOUu6/09is5Lk2CBWZhtzPBKqQnp7P2UfcjCUatJOopsWpzz
6yOEkyV5PZ/VCi2JgOgUiZecU6akcWDg6rfaJSjVf3n5NM9Bl79GCmG9r5jNy/L3D4V0jMwoJoyM
bEWGnST5dj/kZLiib/Eifucz+DgWqShZHM8wklc0CssZsY9XKhOQ2XM5B0GJWlIDIzUJCwuocoAK
5rm9RKYfoUgNXe4WOkJh7XaUdxBsirkvMoWQCrSeyC6Iil4mQ2gMlT2/cvZJSwFlSMNBkloLTWub
fIu9vI7SrOgLL2rf3o0KK8VumM9ELezTkm3p/uinzPL108yC28XBmNu0+Xqw/Bp58/2YJxM4BaVq
8CqZUj0RkVb70/F7kD0M4WAVHuZJlNcy7RW5QO7UUtYsNwJrCTudVAefowexBKdddpPo8+oE6rR5
6P6ANWNjToLw2wnUpv+azXmB8pG3KBnz6pgoIrz30FDynCN7lpOp9Qq0M2hC6f5RktLSS2MuZJ7V
LZUCkFAYuXZwKz7RB0Shfh3xIW3U2m9eq73Rp2y1RuAQeTa+zUpRRiv9lD/I7uLSatiQx8sZ++6x
PKBs2tDJzRS1CoWTa6AstJuWaESO7qn9T6XHMl1jZfCpGUnZcSiQ8a0qxPxffNclIGPZgtWI/fNM
Vcb3mma0vMz/Aa5PSxCKHCIexS9rObNO5VUuOh1uTwIOkheF1CK3KJSOwkycI9s/2wIgcdBZwd5F
OerC8PahxF4jtcrWzc2BO2DtrnKiOAZMyz5kCqY/OtPjVxXazoaNzEOOGm96Zsy3/XvMBn2pV87a
9itVIDwTQh+J/Cf6JIVM+2sHjVes0eJlcxTu4aH+qyerFhBwytUPcJbtGXaEZy/RkQ3qGE0dRIPU
wwu7s0+AlkARlo0hSrbDUjFkKr3c3BQtdm4XsmQa0yHp/Mscx0FFo/mgMsXveGFX7d/8vgg5PQin
mkoL3IkRymecUstjGZ89U0ZoNZQweVu2PqXFzhmDLacovrtYtqnxqghAzxgksXc1qN0N+lPN/fQQ
SY1Ihl1admFlqHDyUMeUbMl45l/61+cNN7AuMbs04tbVuY0QvVChxJw7UQAyhKX1zNOT1B9URTg1
YIUNWAJrKcdz7VKIwZFTr8vn93ClOg5tQUHO3+t1vkM3LcsdRV676+C4GM7Y9uvuiW/SAfOPDetx
MzM8V1QBGyCQR6NFYq+oNm3KIFwnceH88frMg9DQ4MiAOsTccMU7hp/uTQbSE1EPyBFjHQaUEVqQ
Yh1vqwUmbSVEsM1ZoDL4AqUMnvxTp/KUf5YuQvocmuMp+oY+IHoQV6h5+AC37uABvSYYsvz+g8Ri
NldH6fz2YX7z3InWyhKQBHttmRYTo0o/lyxtdnDuDX4jtUhwmGF+1RzxZKLdYo8Cib0q01M3q1K2
bb6o20Zj3VUb4CzGJ1d43x0TnnirYEcoqcgiL/eu46tTDKruQnDIJilT41K9SgQXES7u4npZ0ohw
MN1Zl8Q3YvIRo8SVT+OSRZ0tHOXv8JdyD1kpQYhJntQhmgvx7BzaTJtxG9Ex/mSq9SknnR3G9wpr
ym99iiOMU9IoDXjKfrES7+ehtyJk7+L4VE5a3q1U7Ddq+U33H9S/L+EM2crRuuPIFaZmBijelF1b
k9VbCfxdyB6RLNUFO/tBLN1tXDJKQny+6vp47zscHlU/WA50JYPIDGrMFDvUMTaII6UOct1uoWJk
xXvTg2u2XHg//JboAKxebNN/PlOJ1XalRc55ytIESu+L2O9nee5qHhNpG9qG+BpNdYi/knACCBzv
1YJCEUxYEcKOvsAiX2prqSNYaLAbdNrHztSEgKpG2pOMdCCSgv/Zagsizi61gWstZc1g2DaeBB1z
iVy1T0QcCHuXsTYOJD54MrhnYNK6+TVzprMAJfDeEG3gFftAsRCwKHM5yo14A20ZtyXjpd7lvDXy
ouo2b1KxoWhPNvN6FhRQAorJLpJFdocFJBkahA9+n8lvGxiiSDm7kWT1UX5RIdXkhlZwLBkew68W
IO53Xr4tjrUMWQB9uFAJQGKV083wdD5yeVM+QnOJmE1txKIO6Lq5wgnl7Rd/sa5Fengm+0pJ82O3
JSwN4z0Z6P9d1i/kanuCwTCYFtY/3tqMhSpBd+gYLBZyI1sRlN42zG/+iPUx1dr359KNdWmVKKcR
7HRAr5vZn3yZrIqQgLlIc6a70yMubPnS1PpEGsFjTCxMTAfchwdQcBZpc/0PD7QtxMKIzcBvPhz4
Z8xgdANc42YElrr6NRs7b7hOezzZioKADNHvslaIeYwzZH+/qQf03EmLB24c7Vh5A84p54YM561l
LGHqXl085BoEgaz7FpLgckR295Jy2sZFH98f4GljXectxmSCJmQO9gNL/Bk2rinkXNee0zFaX0ti
CMFjsI8JGKiwHgAccNdYGvh/f1VTqItPbpZnyN83YKz9lekv/DgttzjbIoWnv6SPvObqYEu5FHJd
0D86jD4jeswimcPQwRgOBLNV5g43h3CqYnFyTMeOFTdjHij2piz/k8LW3L7A9YY6qpoprsofsXgV
8IBhWs1noVSCEILL2kvkdnPtlLRwSc2TORe6qQcU4l51tuAVsswbbeOLXnC9ZlCQ9nLt17pQT2pm
N3Em8w1vgeipQpPfi6sr5/hqAgp1fc05epibHIQgnoNdrdYjiapAXbIvXApotpaVmRxLLNqQNR+3
ToPjFUNGPKgVpax86/+HM86juGb2NoU05Xjcm21XBsxfN3a+mLOjgDiym88HwGNGGreY9+7CXkJ/
fRo5VTRS5lW6B0tRUYodRwOdmvf4tfSP+zd7yLvYJKnv3RPL7mGhcz6I2uwoz7I1TZqRvOqgie1/
eR1f8TQhWvef+0RqEzMSiC5OlvXAlCPj8SsL0qejntJZ/Ei5YotW4aLPbPoK+xBHwNDRlysYfCU1
TdMwgr0lA56g24k13DdZ5ePMfSAayE2vcmxMLOP5VUsQjklUVHlsgmSVDI8z6B0FowaD7J+xmFlM
EWYYOBut2DcIhTKATp/FPhx7DOX80++qZoyFg09qZkMIknbZuL6WHUJHsCrCbSIBCfsPOisMYzPt
PhHsNUaVisQxg0DJU5G5EkLN1McJX1+FDC+66ZEnOlRokin8MKuy1V7ohabfWMSOuVurgPzLJBH3
t+cUut5FC1XEC9D+aH9Hk2vGet0Yp+mSVS1nBm1/fEQssniSAd7kKceuvrgiUffERI85hy8yDM05
aHO1j7EAskXxQ1qTDthpqofK8tQEIDFT4sn7K7uHw/tj1aHVFcGkpSy58ZifEB5ULffVBxAav6go
DTeXXYGpukAVGFnr66I0FoYfRB+SeIqVZmm+jUMNqqMPJi9uZse6/vdjrsoAWtRWRaBGxK6DUFxU
4v5UHbBHouNfAVabe7NO10hGroWo2+NqjN9rNOW6MeXNPz0l+FBj8gPyepwXsWfiKF+s1JQTxgnl
ZfdeC2f838tMoYw5QvYpdVLFvlLYZpd8Hwi9Kk8AX8Pokymth4v+34MN6slsBVoMXz/o11oWtkev
k3Y+uneI0+Zhi1ivPRKn9uq8AEp6n0KqT7fg7vXqRT9QAMAMeV9EH/dgErkuDlonUAPMiro5DzOQ
NZnsykvcniAES0USQ9S5hEU+AJKr0G+Kk/x/8QFfyPCk26aDTCsk0dhDh7xUU14MkWjHVoGtXBIw
RaiJB1mP0bJUZSbGXY5F/3UYZ+5A3RAyTh2AeJBpnquc1iwZ9OtFZW42HqmyB511nCukKV86V3Vs
MklSzc8DxbgAU+sZOTxo5oPVFQmOpzaA7uMnxzSiOhTesNDcYacEHoNP45o22TxTY9GUHjHhx8Ic
Am9wJn7wKZQNVYrD01+UASAjcMLOUQ4I8xLqFB6i92xk0yArobzrQGTplOtspDDb2Y32cQfPQ8z/
n1Al4BVcvI66TJZpuIVMg4V4SeaUqc7kEspS0DiWXT4ZSeNlccnFnWu9E9LZ/Fh/k0Mv0A+QUNLb
Dj/u9NfAqAA4j2RhETIWx/bqWdc8WI3S19AP1+yKTLxLQhSp/0J9dSTr8xRtYpEDV2KBreBkwzVw
I+W2//HWkqtsk28NIN8wpqjIPxjKLxyVt6vCm3ntxVqrX47rUk57n2Xr1tM5FJajOxfI35WSf8cq
HInfx5eM5uyFJpjlXLe7AY9cz8qDeVzWa1Z5MA07rHUQSQUMPsc5t4oa+rUrL4Pbu+RiRAC+Mbw/
gUkK0RyRbccKaRFJ5FDX7eKd5gCA7fIUFfeRhlVquCs35f95P3KDQkevIlNj8Idzw6E8IT/5nJAt
yd3j4bDQgUuSRYKymBi6/sN5trsZStJ6you3ptC+kBpdjmzT0xzRX8szfYuvThTKVI1FKOqcHNbS
TKj7tS1fTFRbOew8/mWVNNUAxTVWDCuqBmO8DZ9aBMIAgC3okFGqAaQF5CkHtkkntASUcDufOXPs
jxpRCXyeO/o1nyBvzozPLfPKbGug7o1pjE2zRWRxPMBzX76kYqK+jgm2bPR0sCY+nmOQlBoVMd3E
FfcUpalDBfdak9X67IPZeE+8X8J8uqxBtgknxTS6CNcRtAQx3k7T7ZDIi3+JYFuZ7EyP0dn6KBwD
iRC4ahOJsOhVqiUVyaUdgvTpE/NzHwLViM0cJmcnGmjTvMCH/yL36KJkmKqRyug1FBl6eAqNiVB/
tfYX+A/7cda5fh6p4faWD0XPLGtUApJprxS1b5OrkdTI58swmjImdCR05WqZmpXJuLf+NSUZ128t
8IyQaXRNOWLloIWCXYlxy1QuXW/CZvli95XYzQnesArxkUmY71P+MRi+hY+woTLEWuTF8pnysKds
bTLEbJ4diA/ON4+PYbRijMyWbvix3ZRVK28cGbj4FCuDOD9Tf34W36D2aoBxIP1pu7EfX/8h7rv4
/jjb9sVvPM6Y9sAS87qo+PoWulkNAPhaDpL91rWB3vy7Zn5zzKmzAX0UhOkSVYj9VEF5QVseb25t
AgZMV3HA6Z/fIQ63uYpYnxaBASXZZdPwAt3KlzC/FMelGslyO77Dx5fS08DGRlFnGKjZr9FDtMqz
TgsUEESii6y7SNyycURfWFpgOyJxf/oaACe9l4SzbvZlyC4sS//aYClMObcrEzFq+BcxAvJ8VXs8
jDl8YnT4OQX7+7t7jVRrGXbv3jfoFRfFItOIYPInw0vuMreHCLZt1oaGSFvv7TS75P7CDxs/GL7t
3wa/kT08dP7A1ZnGS8Gkz637x2s37SkRLXVmQSSW0nRpVjNR2Hq7SZbDxHGOE9FqpIy39cSpg0Pb
WaP4oreBBrbO4NKb6yldxO3BjbmqGNN/xuBStokp+P2nhQzNFVtL9sgtjh18OyJhcOAc6127mAWS
zyR9izDT/ejGQNNY6BIar9odLdR2va+tLjZyowJW9wlVrEPfSu8tIcqgfqoRVdcGI5f2xnMa67WY
BV/AgElBSpnAFZQG3RdxIQFFCSkS7tILgR6U8aGgGqVWPNB487ahKvgRq9F02km9Ha2vDLABovXs
NdcQhluqhpzu3RSjjuiwPo+AXU0Q3v7uZ46OzsPMy4rFGl1KzMyAk2dYyO41Fy0/X45t9r34S+R6
nNbwyGSM38biTW4TIPLkDjd4FISD+h53dEH4P8wiJjCAI3Ny1P3WuK8ZdaNcUnKs9UZ0AboCMO6R
SMR5CM2DTJwwSC3qOzxnPAEO5/lUpWqdXupMQ5lff3iB7KyjwtUAnngj3D6YWnOh35aCcQrlqVlz
128zhot8xEDi6/dnkF2pHSwsJpSfyBtWXr/IlT9PVqQvDyebT6AKS0pb9ShEEq9AIbLIKG38/Igf
tGABRhjKCdiRPr717DDcyYllWLS5RIAamCv8c28OjTB6p7xnYpkAU0MLVHrLrrMC/ootVbOcDm2Y
LeWvsz3O7HSnD+ofwW/8Z0r6B1nMZay56giTJ9HoxVjYXO6JSLs/pc9ntGVlsN/uf5FguxcpMuVb
n4wWiUpxgpNek2rkeSq236KamsMI13P9I7WTazMLl4JWK0u1WLQSm++6i844KS5hMHrKVEhkoPQR
vcALLh9HPuOjlvDvuSvcrXVhKxAeF+j491jFvhjwWdIVLnsyB6JFjOLxQTEsmwdYXNSfygqrsBRF
utWGxLujLPrF0vb+IchzWsu88GD2mT1qHQlj/+WW3CxGbxjrv8pfDwabwSvKjNp5lBp41HTrVYwZ
/NP10QjxMpHdffTeCysyFS6Q8jo2kMyrHePhOCrJrN6AVm1PLNtFjMrG2BuI+6kAN8LxShFFtE6P
Oss4MEcEW4FkXaQjvUo+FrzAsgSAk6zqwdFdHcL4vYXs8ESD1ZklDpw/SUFJp+YHKG9sPpE43oXB
g44woQkpn2zjBrZG1OXLG8OZshTGqeOU87RGhcCGN3W1Og0sb2Dl+1zkVuROcdXAe9EEI2+oQgTR
tWyCDKPxLeFxgXSP4gFmuuGaNiScgtIWDLUu+pnPspvmFn5y3GdxffsAojxd8ZrOfIEo2EBYcuj0
4uFqEIFNsnDjm8ynifjO2yTLTF3scd+lFNEQEsFliVEnJSVC6Jg3fiW82WM3ysJ8jVaIbKEY1mpF
NTlsO2swSTGXLUD+QPJPNlKvPOU/w5iCMFCm1d2/SnOEI87cvEjYRtEh2oufjtv21nehg+KA6jRU
UGRwRjtrpYl8fa+9am16T+uvec7oUf6iv9iosMysg5suLoxYQBBU5/+jOcuUZ+YigxNWFJ0+VIpN
kCnQ4qyHjGeD32M1tH/ELpuk0xCI7zoGm88Ut3NU6YrJNpgyTtABm/eeKmoPduGVtMZxpq3wvdqh
whnDh/XzbO2fkitLCwkuzbP4Eluy/yv/fTLdkntIQCkoKMtmjggggNwxZ8HwsNSzcMLJsH3HOHci
aAtzHyWQsH08y2KPCqIzPyXAoXNyV8SQ+4a3E7xwErvYHjovzuxXH8h3iu4FTpHSFjnRh1HTOlL3
Sku4scwCrv047VBIOBYKN1KDsB4qrtRgoZ5E+6VmM5DkviHGzIIOkrj7ItOb0Jbbb0KIHWN8gBBr
126qtPYIzbvVueMPuiH5Fmz6NMX3FVRmRo/ngHWRo0SNjss0GCL+tkl3g0K3NTtv23tWJgaZNyG0
4IJbtZIXURVzRB5ATPMifJIOQjLkFO1CZXVv8xOSETtGicWvwgYrVcLsigeIaqYfK1jDbJ3qYB/I
fZNEE9FI4lmCOc0StXP22zHj7mmqMZZ9M9x8w1T9/kMtvgOE9Xw6axVJb6Dbl5q82l+Pj0qG2rgj
uXf4nis6n5WRz489bAaByHG1iui5xmVM6O72BbAfxjUkUozJL0Nv0RbV6wOJkeJJJ8UFttNmXBDt
Hse5WT0M20EDRw+HzrC/uuGJlMRZk02byWjkGD40/H0/acknKz7JxqukQDZgEdGlXa5Ls4FbzE91
mDbX8QBB6G7qG/7iG4I9C/ViPTSdULGXV+1ArkBHliFnnxMU9EqunTdI4zoTU82oIvwAOcs7+z/E
ROzjJw9FDjmMidI6MM+3blxgHLF5loJ91td2tFbZV0gADrxZHRrsQnpb82lk7Teba4Wb1SrLBT6b
/chNTK8xjIHYauiQXr7ZX+TOf92yyOL0qe/0/2Aj1fu+Iar4lkzKdVIq3rDLROBkOfUt5GxoBB9w
rcsBKzg+s1T3XZokcjdN0LQ7qrm+AJBqiyqWHv8lWjTswgTy+eP4cxMGEM51fBVheYXWkOUeWwXe
RsgzYnB6PEM64qSlsWeKnyybZ8SaNLYlBfS0BvjJALpPq7wzuO+vS/IWUckhp20vgF23HjMmSOYj
C/2h7J/fWbV6ukkVB47dMrCmYEyBJa+QGbnCMfLHi5mJLcoihS3u1XsyWpCbqi0wNCRfAELSovCZ
IDlzOuc6fnT2mxa+b6utJMJAhiYHU9VdwO1UvhqNGnOe05iiGVNL9DAkDbfIof9OFIswleS/CK4w
W4ES52RDs+uxi22FG/ygdPDC9oJEA+PasBoM2w7XvN5zTQRdBme9EJY3dhWgFAsauT/Pydm/9RBI
wyEvnfb3F+yivA0a9OVMmbpMX0hJ6Xr/MWwF3lH3/jwt6uBsotRtULps94yxLKPJNh+XLoYtJJRi
GPwQ5Jak90qQUvmkmdxS5sNO3y5UHxXrr8uf6aElWN2rkZUnuJxbSETaVU0N22xkjaQfBrnxcmTY
8j+duCIq6u1FS0uQrEFf+M+3BEL84IsyaLsUJg02Cyz3UOD8rKIDV7ZM+Q9R5VXG42UofO7WfRqM
ashdQ9LahCxPjZaVbLRZ+F51+UnTwnscdAWyeSmdVBeKxlsrWYA9VNFbZ+c+ShcOM4exMQse+53y
N6T3Z6J+6A88kyT3Qv/CGIcGp/mQdTgnAZsob9BJWTYwvE8Nh5TRPzRbDFMVq0CsHHOdjvSCYqML
Z8Ukq7T6bKND0K7cyY6owCen4BQfgRqujSFtrnWrR1d9VtPhZNqWWFmM1oGKGjNL3XOmpF28LLtA
P8vqtYRYMFNAArzY8PO5oVaiWNi6BxKZPnW4V3FwBwqcD8rRsDZYuirj8W+zs5de2t9ZIlDd3S8l
u8iB4Douqinaw/2p7MFAd7Buyxh3lJdUHhDXZWn6JenvqzlP1rY5wzxdDffmoGPNqSEDitQZIwzv
6VBgwkShepF3ywvH6RG+i6vLhKcySzBA3iQWWNH0v+LFM+vTi6GQNKOeZcUZOJWC+X/q7lm/TGMT
xPki3OofwygHuxdXhzyJp/z0dbkeSXSsRscZ31PquCijejaNm9weeCdXWzDwpPsMrQEaNIQtNA/d
sIKQtkgeUaS7yqalpOfYeeulMG/ewBKUEQ4hp+C36xUS9arsOKDbDrl+cwGTRUEokYWRJDD4rxbm
Oa30LtTx7KThbgBJ5W5yeMXMWpQe4kEBzbxpBP2LMR1eNrMTwS4K90FVw75HFFRU7ZDStTGvmsLC
j9eyK6HgeOORjLuptJoAMSAsJ0huIDWMUDx9/ArPEwbrGCoSAFgN3x9jk3tVKlGSdbgweB7sTKxj
uj9fYpOgdihsPsc9lS385ZpvchjYAuO0kiUFVH+EqfkdG+Mam9HyDYjMLrk1GEW/AumhkII5ZXxo
tx96LTgUvtefRvv52lWAli8XiZsKyOUbEwpM0w1Isns6Jduydmq0kJ+mhG50ZE1YiQKenukIGawP
FX24H0FWVbqSiOuTTeH57EaUeqi2o+jK0Zt/Qy+0KzrMDg0fa1hy7gvlSfbh0jOhtYmhj6NWyaBj
fk5aUEYcP9YRtw1T7JB2lq6BlOwq9WFXO7QBXT/GlTvrMibCg6m84KldzRB3LZi+Tg93JDR5C/4r
zOWyEamxK4SCiTdM7nTmm1v7XrUGq2/y1lxsfxEENqikB3kTYGEYHzTV3aAWelC8paw/OcMNYGDW
DLrlZ2f0jCp5EESoYyULMy7BkpivZjOjHwz4ix8HVx42U6Kq3QgXqzhpcr7d2O3WM7eZd1Lxt7DG
pQvgcgMSV8ZQaUf6s+8hwPXSVlQGYRlt+6CprVKUR0w/jrWuBe1Mue1C6G4BGD1i/oX2et2Gq27z
hk9UlY4G2xJVUGQqAnrEDKNazGKx3wOji934N7qoKpREe7s7U3tX2R2QpyWvHIWZQB/zWSwOucdp
K/UCtq6z2YNNdks9Hk6WcOQYRKqyI3Q4nDsNXu888zPve/o1aHtkb+9XOIlVQq5JJsCOzQLmLard
pXp04DxY6PPP1uC0YON5a2e6/5rfU6y20csVj5AW+2TDuBoe6gYK46lgQhRzbfd7RIxPcUEykVXs
S9PYC1msHC1wyOu9I+7fq1vCVgMgnhRHtPq2/L5JqacxKZo5Me+aJsLE4AbphRUrtQgA43AaqRKa
YZMlIFwd6Zjmw5j0vcVj0UYUgnNoNaTKZBLohQGGDHDr0/RzTw5lrV7bNUAF/Zzxrdj47fQqdMS/
jNVvr7lPdpwBCz+xZlPS3Tog5imGqdnW7Fhymef4mebJ1xflxmUtVGevvohJS1SutsGgoMnY5j+E
xMcFlZO3YuXTXKxE597n6m5M9bDnpPbiUjpFo8OQhMWATFGkBYTyleXQedFDRJQhxsaKKCrPB7ze
rCdc5PvxyyxsXYpHTsIfIagQZnTTuSYV84X6AlI3++9uiGYXRttlTVrWhpU1gmAf2EMqSkE0Vq0v
q4/Gxtf98pMGH+LML+/YNpZiDVrrCn1mGY3zBx6VlyvCmnHN1+/2i78K0vmGE1FSjrPnC6LEoD7O
s4XRcDieHFHzDExRw0zmDF81Aaf2PKodUYxGxZbAocwXNoDX2diLodqTFuFbUnq0uLaY842/ejOS
Su3D7unzkQibEdwAopSmg8+i+QctrvWi2wO32T/9nl714xeKv2t2NGE87rI5jGcuO+UqdJ4YR79N
XiFJBDM5hHOxAoQJhqcUfPeCFSanNjzgMgJz+jDYKfAvWD/82N50nHfs4Q0JZRThVzlZIlOWHMHo
aPck8Ir/6CaVuOlA+Ty4COtjbq2Rmou5JgTVMhpfylbPxTb0NUBkWg/0Sy8gx24U1RJWSFexpizE
POohU4AQi1N+M5OqBXESnRAsW+P9Haykoi89tbcnsLux10YBytNcs2NW6sb6f5od3LYql8c5KREO
Hhmbk6yZiRCa6PUtFABxO5kOLAMqgV/uFkZt+HIpSiweRauihZj/I0qDkyBPFmBv1/7Ye6gXo2ne
0FUF05YYlWC4miyI/6PGf7TIJhk/M1eYu6bWUf9UWoJl1/JSdn2545UufAQZSEt6ZtCpDQDAV+lM
ffzo6+bByTRof0s95ScjrKujJ7VIlDicL0kZ+t4+bIP7Ui+BoBniDYIRQ3fT+T2aE2XoQ4iOX1HZ
SFI1mMa0WGBlMKGKU31BggUb+fUgMKMpbXFAgk373x9B5drCMlA/RFuaszswvSBiOLw3xDoBBFnf
xB9uTKZr4ek6YJanD9uLxxTlU2CsYf3yvxR0ApQS4qt6ll6G5/mWULkQC+Ps8pR/UhlekhmzKseT
/dWIE0p9/HBuqjoTGOLJypwtoklNIgfBQne4uE27oKfg8BNKp4p7TfIrQLa7CAbXosyGOOQJhwIl
Bxco1DGmhQGxzGfpve6ME4bMNfTCxkJqwzCn/J5XaNbbPxyMvDwpADeFgJyqIFQr9kT2UhWRubzk
1xyWA04at1aE2WEDa9W+71V+bTCil8KVKYGhehLVZ/3DftujF4LRhg1bWqHhmnMs2pjwVXbKrd1F
fXMkYD1w8nnd6PHBetaBUq519snqSEtG0G+hV8v688KFZGfzLtTPneoTLb9pvXDh6bTFDoAeye3n
KoqDeBUBasADxAcQrRpx+12B3IWAqkzCMmsDnrRqp4ByhRKdQXRwZWXtwR9zLPLUc5pdRPUTvndu
OojDRPZ+C8hRU37Iiqjo19DgRjcsJjJ9wVI02JioGW1FdWqOdDZImPw6gOaKrQvuonELO5mPiVMz
MVKn4YBGUYntIf4qHpJDuwTxvZ/okbVDiLjAU3u6FUDqD5XBsvUAzuwTWptNWdVjqPt9W1OnQgVj
lgrrYDGWkDJP7NgMgMwj9ZV5QrNhV5Xr+TAkloKZk9dJu+WEXNF9gkZizV2BvhV0+ZzvLNcZ9R2a
iYDNy0uBBaqyiL+8Gc40xzooA2B6pyO4lZcdxnZ+IF1TpYZ0+htF9aAcHZm2xKFCw92BdvJVQIlj
bCu1FT9GRfvfWp5wejbcs2NXIIYeDmkollJLjoAJk/KNhB0FqAEExUctT4JzLTJqTWrWVoZ4lux9
GctJUFF1bIinADOi32jDIylL/ueRnNa2s/cahWAA5JiKZqY32GoQHNjS1qxLzuEW1zjKeg18W5br
q9sbbzokdNUzopZBnEBVcrsJuf/zLl6frP9yeOlElVMi1sV9mAtSXe1m/96nE3Rx/GzmrbMUUKWK
+sn7sAPYmSsuwIb8H5DvQjBBNreJkmgpHjnIuE5ck7b6YPrJtrTLKJ0SwakUB9vL86JM66XQR5S3
ODW7PgfTFvGoumUo/f40giPvkmbvG3Wvva0ScD8La4PqxH+df1oPj4JkLCL2pOLB3iXUJPePPl7E
/jCeFwVME3xrTf70wiEwd6jmUdKLrnLAPatytzSn1d6sQczLR+ABiilKbk0mlzcjJ6OxGXjXz1bh
/HkmouzUlgrOHftWQVcfitOlsEbmgTevaxBbH+B+JBlpO51tm3497Cy0lR9BDPvfzSL18xWBhxNj
AeIZP6LdiboXG2ygtAA3/edeKZdCX7muFyOUANVAEm7gv+5EYjZhJrxJsQMrDRSGhaIR9hFGYAmU
yAL79hjaxGAyTIJtY8tp0Z5AHG5XYPF6gKES6OP2eHKoUNqceVa2kLutR5+HMArdFlXy+Bvg4hVL
br68hGBItQ9EX+3i1fRJ8s5mgXStmNSPPSylO+o0mB3ppGdwGY1RsvryF1Lu/sEzMAYfY1EAyGRC
+o9YLmfg5r06NrH5CNR7ycna2uJJI3yDjtlqou4JM2/vJw/zeQzPe6j0BtOOg1JoGtksyKOTUtLN
9HVcPmklV37H4aA1kGwh9cW8jc8DfRTXJrsRP23qiJJKG+XKbCogsBgbQ99J5CdytpljqQZqRLFy
lrArVKKY5A8dzM3Nkx8fEoHbKx3iXtdV6Zcnp/qtY3A1c99eTg0AGWLgNYIkiRKv5Mk5/LN/OFrD
1JRGUzyjlc4LbYFaYijSTJqfmN0WmWkWkg6utAhM8OUNyX7Izyp4Kfw+FPUX0yaZUI4e1nrKQ5Ei
2jFSCv35kwRyWizfo5R4cPZoMvGB7p0N79I1+O9r0YXEtUjU4cUGf9FALq56sDCzZ0kyMW26mG4q
9pTRs9It6rHfo20QhY10ZR6s3bfj1auLCIuA3cu2xIaTy07V+s/iXYeP1H9Dsz3SLb28oZCRtd78
kADj7K0FKTvQaqN9NvJ11LvkLBrhOVvd3gI5zRL1klWMvGus81Vdpj5SDtRmDByHBMaJ4I2knwEf
NECpLU/DoT756rZIVuTz9VDem3gk277cTqnmoGqVeYPH/Cjo4cbeihjxYOa8nCHzTx+Znurji44a
tCsJPl25g0bzcv90b7NZNmi+2HEsLVi/Hw3H1H88+24cjn0W5zOVnYKkU3Rqw4ZmH8yJRguWFPFW
h2XYYv7+/+dpYytcBooxyttlbmomfti6rhUz6pj5Y9laemhaZCys8qpog4whYQtxqmISGxrpvp/q
8Y6ItVbRRfzEPliv2aR15+vWMOvdeYu6jM611rIMag9rTPLD+TQJfXbfH+tCIlB43ZJpYCpYOQg1
QYYUbXjWd8EN/0D1M+EJcRtTUwMPeU6qXEDwlPXW3GDRel7SmNxSREbhe8o7cFH8jtpLZK1Nypoq
x2UT+cwSTV9FyUpM3K7nLyx5lmHctBGZNW5DhAAP5j06KBZbvrqUnIdRyvGdFFRoN5geI0X0rQhU
cPZC5gUh1x7XqlvCvNx+zIbzetnt/7vlY0wuqlcrEePEncw5uGlb5o/7mqm01JOOzoPNuXzorPZ1
7KX5lsJmFyvXyk7tLqEB6DIrnSUdurA8STXcTLqO5R2al9IhWP3OtCwO9UFsjcLHyzld1RmfwUAp
caEtXEagWIN1snjGbyGJyB+YAqDgW8y2O6asW2ChqQUjPiSW/7NtBEMbG/CNfU7hFtPlOTAuIvmp
2qGUk2ura7ifno96TQJmBdmnFTgyOvvz1p2iRJkaGMY+TCCS/k9SFwuWDOhMK01zzyCVCn+qt82U
VKIRiWNWdXhZ78Z5ln1FL82iaAWSn8gSxc2LdUpx9g1C3E9mlP9bgThuJCUD+sDgZ0VqZ/MRHDuv
NFN2QayLA/rX+5AO7PhKQLjAeD3wKiyHM16gQ4PL4AccBwM/jqrZTqoGJix6hcQ7s2vLZSoooUZU
B+CBjo96q0cz9NFjcs9oD0eVG/l39gJFPor+levnsTXDoroFvlYpPtIL/9GnKrnNTwD/Kd/ftHTe
RaR46l8yCz/MXcdnaUX36ZEdVdRv6GoHRKJu1VXZIXUspwr5dyzRj2iurfSWiHWDdDlEMfYjW1ha
Vq2K5kvRNllZRfDEoj4DnkKM1oS9S5aGo2FmqWYOpbpfwLPqzEyGMfCna55NPBq9tUd7PVo01G9i
G3WbFWL8343KhKSGVHVZQaR7hkIaR3zTVhs2yYkkgOZSgK6O9cuuQ5taMZmdn2vSDHIU6ctQCREK
S3ISVpiaEKnoqSbQckyVewOdAFk9wKMBkT9uYhbSi93qBlV337CwyXJcq7JqoMTUGN0QvdQibJHw
UQ6TOlRQX5Rwams7v+WVfjKwUZgjtMDCShj2JF2JDh5CVjbHfq27wxSlVVAXjM4XtDY46C0eep7a
ut9LHpM7X9Dn7pKKWO6DoRhD0X7NUGySpcdRRAh2DuAODHWOX21nb2U+MIlPiLwsrMvUZ1LtiJ5u
gqx+u2I5sWFtHhitVLurR3VaP8MFSxHIhF3IWlsZI4WlB/yXL4cgmJv2dGZgbcIvFBs3gDHEJqnh
jc7ciwYpSoo7fCa91jq2AYXqcGCwGJmgKGJ3v/P+WQR3eaAa45zBeIPwceYuCSOHtzZC/JDM5cO9
90cGeAkjR0LfpwBdEXx1IW52tIWANEMKunCMIxG7QHYo31PPE1ZQkpadxZDzJeoy812ugVoJDgMC
tRP9HYMa+BiDa7Hb2vlnmMxuJvgQlrmqIBdoIzhM2yD/2RE+dk3EuVAvomDaAYxjGh+GkyU1WDB2
bgdPCwusq1ioIYP38B+pHAXn8H9VoCX13yZhaCVk/i5bKW9M9+5TF6mpEWi+mD99wOEAJuimlJrv
L5F8KPJEwQUgScJ5ZURNty3/ASD9+ezaa4XXZe6g+Kmca4Nw0fu7kwRO8NxO/nKFMbimsHQ6n78Y
sm4chqQveq9Zpmsnw+wP61TvjUjOnAcnrICtyImDsEISelE2DBCwGqHz9xhvJhtoFZXYUhQCP/aE
4BO7B0q6Jd601Lv8jhWv7XZqSSxBIP3eDnwAd0q588iNyCCNTX65EDVfBD7Bn6IytMxWt+08rlqb
1cM+ZlMzmLQuCOrSfQ46DJW5C2EOk5/ETzqKCJ8YXvQ8WPrXe4aLT4aKlH1owAwI9FWe2S81Ha7q
VpgIP1NJ1jOGp3BxfNpoEEpl7ERpCP6XBQwmt2FxiEjs7mEjFA99YqwjD+Z6PnPF6DxOaA4vakvL
V9UdakJDjM7yMjzQl9TNCggL84MMx9q+dRBQD8162zQpz8rCHkWbCSMrv83HimAKFX5uRyxiGx/C
PZTVGYe/T6KmZp9mTHeJonB7WyY3dWLdIp7UP2LAmqW99fPS6kNO3gbnw31bWvwV4wkdek6MXtsR
pi/kSs/J6vpDBx44I1TNxU1FC83qkbJR5BJTs1OUfCl6Uxfnlafhfia5xdIUsTs3mCDO8Kio78QU
h6oYdbJ4HLOC9XctXaUYK3wku19PkzVglK2LCpOLG99pqswEmPm89vsLvVrB7DoJWvbRP8soSi+z
ZJmzbaD7KguxHM/4QxPBpOjJGFmSLS0ZvfngdHdu6CnveLKlxn659U1GLG76X4/0o5slskVm3qZb
sEMw5mzTLVo48+x7zka+jzDSgGeNGd1STEIONu4JIbxTImr6dcy0zeX89UB3lD4BmVAeU2nXl5qu
oimwMGzSFWXFlOf+7oqPnR56Mv2g2rHEP6GjY3wPoonqId5hv31zVP1z8ykVVPW6rBv4OjllvHvs
Pk0ImuwW364aPiSXHtWmef9CTlfmPTOew0qjctzBDnwQRY3Fb+pqC4yqWqX+jIGdje1QPL5eHEhN
Ns0Fdl+Iinw9ik6+Gqu0myvlBtpq3IMLHDd0Gc1q2w4ypPZ1ypez6hGX5Yr8n3bO/b5uSpylp8Wd
NDqOxFf4qh5D3Sv9+YxZZBDJetludnalddT+DVCv9rW4kjDC/jW43aXf8XbkNRxCr203ywxCLyZZ
QbN0wfA0NKIkOcB1J8tPjJqK/HLW6/SRu3aZWeAbrrceHx+MWKErmfRPJdSx28CLTiA+TjZVrfmb
kjcae1dBzimTVfpy/vWCCFgBZuwzilC/pSKDoeEhkWW68RDWaXIi6GULK2yyKlPHdXsKrCW/QQCq
tl5xmsSS67pw6iwhSDdRJzjk8iO9SOhp1QBBy9NMjEh8w42c92a7JI77VNE6lY4IrE808SlzLOAQ
YOwyn/coAsFWUIj0qBdDWqHGIBXxR29FbjNHWufztL+mxkTvwb4bYCAZ9b4jBLgNG6r4ECE6Wh2J
GooXtbMhB2HEdigios4279abYuGZyCienEfMjOmKbPcmBQnNaY7QaKsfvNF30Iubi+8zwEDmdc+y
R3Ap7NNbA0busfxVmLE6sbnaiieASSGGXk6VNp9sTNYIlRNh2tu5CqC/Wl3O+R2wftr+R1NFlNZm
tebR33RT2Qefhh8eJleyChcOUEzQ0dts9zqASz3lI7IJq6cE68zzD3oiVPIyKsrIoboFAunyDOFS
6M363WUpNo3fVBNBLtUwuxtxraDtNVJmJ8b3tOu4zhKgR2w6qpsG9cUD7a2vorTlSJlWrOCZiB3P
A9V7nis/lpuwPe/ZMzpQw7zywPRkxbLBVKaXPj/WK2ekSl3l1CihqZsujEnXzW+VYv1P3Lm9hAmw
/QLP+cQqMc1dXp7aP/rsR6O+X7mf0DfJbjZJ2P9THQuViaL0dVYTTew6OGHHBZ75v56ikeBO3Azb
rw1Dxac3kwdp/roFWdCAVRZV91AuUXgQZKh9PG4ykFd6VkKS9W4AO5KcCSIpnD9AJpgYFOLataXB
xwFnbLfW/73kFlBvnh/F/Ha5SAOgghmOqEe13O9RFPNzMraWtoYp6KEOCgf73n+xDCO7Kx7U3aor
9We78IT2Ac22Iz0ut4lKc0FjHNLJvqi6fBjOWRh1UvMTverSujEFce9ArVV4W0jjc1f+yHCv0khS
lP27ifDgWztlUvoPEKhCkg40H4ljcps8/1x+he1jbY+1tGjtI3ena6b3MnuFXY9JVMYSEKarxJdH
oIj8KL07WMO4avlROsPXVZlpNnqvHxv0zVyKICBw+mhPmwgRYxix1uxJs0OFiYTMC7d6G7MQ/yCW
iESXr55Jh+zJ+RTgfuoY5kdUFxiZEg+Uj5Uy8W9jWlSHIZNnhTje3DRh7UM52aKQxcq6qdjWrdTc
AnuEIGzsxAM3fGqKzhJQgrVC6P2bfmCFy7+Wt4tj2bvffHVpJLeCbGpgXDH45gFMqfzW+DBjHcgT
NqPyzOXZyE8Fn3gMZ3COZ1g3ouGYvuPL2g4xMYkbgge8m73HCevFBaXDqNuFuZDAgwGoPnghMlkO
+T2KiAfsV7dcso4Mv/BUIOsCGH5nbUGxq3sX10J/Q1ScZRxJRh3K/Gp1LYPJYHqXXCrLxff6JdX9
uEmKfRDs+PZsYgXs9uD9sTBOAcLX+5a1pWmPwSRLxh6CThihy3aOYC6+JnBlA5THpO8DPxDTIIjL
Q6GLE6GAMLJ8PuCHR2K6nFla3y7tPGKosEJx0havkl7AC9HgD3c/hdBmZJErKYkvd28O+VXZlTXO
+kkC4f04izTyyOUUWvCXCIXG50YMjPuwN+St+9LEWUbgzTMDADXjyDFfu2yGs7bTf2MXBNJjk3oW
vU45BZkrmNa4AjIA8IkUQ4qZBUE2WL8pJMTwbFZ+nOB2U79EMVJoYFLSkNNm8oBn4cKgWLr0J5l/
AL+uV9zYuuNZYE8IHCwcg/Ly8ItfB6UK/KAZYZcWUHx84fyY1d1c0aBOpmNmJUsLZQSH1elEo6PZ
c4KFdOgQCANwZ8e1yvnWnmyXO66i/akH9UUVp1owVWuxmcvvp1Y/qvlgdfwzLHxTgPlG9qVP9M7e
p62V5Q+DIpQ/SLSzkQohV8ZntNR8N4Gr+ENazX7ZMtbA39RTKNGP6fYmTUWMi09K0j7vRC6rdMk3
zA85xLZZKf/34zYqehv4HvDKRfGPScUd+Z4DxmZUDP7suqLs8KHXDDqsSNJPJQXx/0Cbn+5qK/Pf
4wr4EF3DiYP4Y95SJO6W6QPjFvQj/yatKBn5C54dqntv14+ZnjAKZh8XRNOV+snShnnxnbGpWVKJ
nQDsyQoUF0nXeKJAvL+1MapdOwuwZbH/pFxJrqVqGUE4osfKamrYXP9M61CZuh5LQO2PC8vkRtcg
kXA4++nTBxhgrV1cEaiiaUuREXE26BgfYq8q2vJQhu7icGx6ykCFub6O/uNGuIgHna6uPaeMGCmS
REalzA2wHgzln7idrndzKiGm/+BkwwnHU/JTcRrBVKVfDLiuQezQUnIg86KqfbvrjgQJhsouaOdi
FO2mjT9FbM870QeVZ/mYcql3bEiFMaRTxwAkOTtVQcIs0lW9qzkwAV6YAGpPkbgAJhwdTDzQ+3Wn
fRQPig9+tKxWS1l81yVYm6qhapPwfu67HPtgl+hqccepIcsR2+4p7h2yhpgXd3KbsfG1HKNU2rGz
BQ9++oiuAn1feUrs0rGE+wc8v8jl2vxhXGjfUxmVemZrzEE7qe81II7nbzT3Xqdyi3yTp6zNcROM
o+DtF6P4N51Qz/DuaTcLdreEiCXadjcp5B2lpGe6jStgOjhGCV3s0eUL+Zl1+/9mFwtI0zveVLQY
Q6PdHwf3ZuX+8dwafzkEKAzHZt8DBUQ3eDtBOFMxittARreKBNv0CNZbMl3Us5vBJaD9hRORytjP
Puw2UkNQhY/czOXeuOVzV3ncPascwobIKoqrhbcoJcYkrAU9eKLV28uZWSFU33YxpCmWPJ5FuSjK
h+S6Hq7VZX1oviJDtsSXYWGbCHQyjbmA3y+OiHhcvwyMe2BuXIS3GGu3GOSceSNEmH94q+qGXdhb
hcxQVq+Xx/b+4RRgAUvSyR0/2WNt3vhmgUFrEnhcnkDv5s+78DbNOoodxiDxjD1RzwSV8Q4nJ0AR
GDSqMOqVcmF9CMOzuDdrFguqT2iT/zGsw/6YeAdCKAArakZepUcoVtwEpy9T7Ib2zwWSSlWwtLRA
FsedBo3W1mLt0QFgdbRltqNtwueS/8aDLRfcIio+VVYi55ITLgoVfEd+ukYAEv8ykxy/C01xVLO8
K4lgj7czYDROgBXHkj9XRTYJV6MefZzv8ooc9MrrakKNBspsmz1oWRyWHYTFkl2cELxC35BoOf27
7dqaurXmbez2T2yPl5nSHxSYt7o6QilZqYItfn0nOj6f2Oox78kvwEwrG8mYS8V/ZpPD13G7nlH4
B2NH6YmqzpvaWgG0yoBMOx7omPQtSuQWav6v4pyPXfGaJPCsbYytCH4Czw7pELMgtRcPaWWSRyW8
h5cDUG6oXFtolRF4KgRCArVHWw8bcsZ84vDSzLWzYvfLzVVtVQmbWO4f0DiYKf6To9XjFH0MSwOK
HNVXKStljHOv2fOSimx7YqkhAMS4d343Twhu8tfPoY7dYF9woLH+S533sfp/H80uzdHio9lLATAx
80dZ8g59dDBAWMYFk9/jwWv4T/Uy8dfh/f9gTDHVbz8kCys2qZrcS2tS32fnyFDcRdg077xSBbrk
OQ+AyxrfvqjInfMMPqWd28auMn4NR0mG12oZu+jBAFLmcaCG+oepjxaxcwlWf/cvcRzl8CCvfUNX
mFSESSoQVXAaDyNteONjIvw92jsZc0/uDQk+VgJGBTForbQDJl0QyggwLHnEBhO0vS+gyd+Nuq8r
rt8jhJhYlfk5REiRfGzbsGkyUNrfYZbL4H8yKs94gCaWWO7qs9rtSsVqKK5Q/AjXFQdafmkVONXb
3IGuKCuhIHsDWudFqeoLxFdhSXvHjYtXBMYc/JCnwJVfHAVTFqQK1CE9rpUemQSereG90stETkEE
AZe4vyNJV9hHYHdN88l7tKth1GYbH02dxauf5Sl0Y690NXIQ81D6Go1sBRWLoWFRs8bpzVmaElOJ
0AAiar/77TOa39nOgxuC9L7lzKW2ZsM2yMSuzvJHd2KAUfuWKBKGM9T2Ti65+lo8QwxVKXeXSPKR
psYaQP+aITwPjofXdAffKxywSipew8SZe2JGAgdOyB8LjNatnfpH2YQvrXXaHLanLLcBRCLho8M8
zi+51GjkZ8jNi93TGy1JqsNt+VDPYjWgfYgIdpxD9ELT5K+BHuAxs3mOtqnX2l1tUMBkM3nkBAQa
LCkpyvyU2Cl9VbkRATC6ktjbA8QXO0k5z4UvMu9C7KEeqtwbBvdVYexlbyiGjQTJUdHQJd1m5Xqs
c3sakZdxz+plgaNv2sSbJ7EKBpByZ1OaSoaazly/q31KF1MQgDbLAV9K28TVWh7hlbMF1T2o/guq
Ska2RqRF0rUOmcdQD4v60p2klN8aBRzPBPF5jM8u6aLmNfsIHNvjNXWcwmTaT5XDISXCf3S2jINQ
zlv1kLrLyjfxHAyKVF39OOQJA0Fa6tDhkGH8gmIPrvqhER11Fvy3tLAeLESgYKiyGBYd4+HrPE4s
7/wzz14l6NXSFrn3ps0C8Kej9gFUR1S1A3P6UbnLUAg7kvg1Sw6v3424V8CHwSpW4uGIYMSO8H3n
UMFc8P1nx95gpD4fzOhzCtTjzBTnVhOshcw6MElBSt9YmrvTXzBhef0iYv6sfhO+5dxCEAmqYqNo
adob5tDA1jRGJNt9Qm69mB5pYSp+KYiTchrCUq+Hiwn0O8SSyWtspBfp/FNYjLCBbocPRz8m45PB
LG+ehGn/XLDK1bQ1JznJv4H7K/RtcGu04aV3oxSsvhX7bRVkYkfqCwRkgSUavqBHacf821MTtADf
z7vTSKWbv14mxiW3XLNyQDylvbHFjaUX6h6DQraV5MMZC2OGQPNEGno0/KzL0rZBmjdQ57xNyCHe
b4Rrj1vXrbpyP3jbmvCaIORh/UDVo2TN63mo2WyXBFrrhqcxMcZ8BvOcGt8WMCykuA0dhEYM9Yp4
OxXc3UbqRZZxpAS71M9Z8elWQnrntaHzKehWwZCbNN8dDCPX+rTRWxFmwH4YCmpiyUd9GAmWNpYh
bSeI6kIWfn0tTn0GgRXSilNdS7BBFuwf3WLz9osLyzTKDvc67uNnaV8+KMTj/a9m3UfSGsHhZvCq
Yd21DdseMePDVToOZ4WhmDC/985OcSxLYc2FRMhRhJE48csqN993j/I0yBlMm3UPfU0C0tC7y0KF
LcNFIgUz1fHz6++SkiudCWB+IkQFpL6Q++tZCdIc5Vsf+/l/I7bVEMfXoABFFUIlymCHzkYtx1kw
WT5j+tVKtjTK7XV7Z7G6Y0ymV5dsCxCenXxpvT8qA7KydQcJNLSiFqxqsd1KlABAoTkdyriPILNN
nOrC0s4VFl9HCmDDnnUzp4NaOBEyucJOtAJDG7HC97xxGltij6dy1rjWYqfgo0tsHYJRXBkJNZhK
iEjQfrgjO6r0dun41HRDxtUwoHrWfhT652PzNaeTN/QYGwehEE092UjRIyuuzwieszBHVEwWtXbp
XOqrnIOa2lV01UPoN4RzG7nvZhJjnzjhpnOXQp5+FO/i9gpPQ51HlkaX9QaMS7cYi8K+z6z2WnfX
tjKvdIFgREaFy007EShXYHQ4HtsqNx5ePH0Ncai12sgNnWuW4ZRVvAnxpsxEpsPHP0dPCkLu8HNJ
aEceEDwo9iIbccyzYOOvJ96kOrUAJrCYty6ZBfpepZANW78y0x1JITXSRLsC/whD3eIu3LhKXgNL
ZSu2GS33bOk1IZrefBDeKz9+5adWA+8UcJz4gbyYUp09sDTtPP6QU+jW985gjogmPa7MySnTcPeZ
yWyx44FPkE1GylM8qnZg+hIg5OQ+2f6j5IkJSKq3o8VeJ9jRskkUmcHYIAuXsY4egnGVYEFjX8Vk
4Ezz2pJAy48YWFHRk1MeZ2jYEAIz8OBbqb1EeLqHAHfVjWgiETK73YFWztUuC6DaV+4hQqDJaJKu
MFugmYKvtyaCAlHuvzpH9NlNAhrWZTFuZme6sQSqLfd+PhA5NQUbxoeqwC/yXTbDJ73peKR7sT6x
9k6lx1KyI28Fv3wfAPUWnfdvQdjy3pMgHSlHt9iaPFniJzSJdcC0lG2Jo1hdn10ruRGjXEi5uASv
kAyLK4rCCLB17DPEubTLc6E6yrt+lURwRo/qCKWXKuWJJt5asSFlpn+bRZSwmd92IQ6WWUoUCkNq
v4zCrZWS/kJY6abiVZevau8NQ87gFlzHfgkq/UpIAtqJciqeh9Fmyj0NwpI0xRY9+WxXrSIg4xPp
8nHGnl3IXZ3dbqeU7lp2cAZzS8KMQMPmH4uzwprV3IUsyMc079Esoh0JzUZ5PnaC8g1/28mtvRwP
Vn8t/+iArRHhAAkeL13IE6AsZ2twLWf8UD+7Vt3RJG1hGEftAVsvm89czmIRuww4YTROsg8nIxHO
0eOomAeaAd4HHDobxijYwtmUvar0iIU7F5CV2C3WDZ8FIo70GdIDaWIaRfhZx3wQsxe7WRfZEfoX
fCeuilGM4SIzKzDD4Oz9Q96WPANhsq2rCBTlxvoaSaeSXWBARABwFrbVQneb4FoNZeaazgHjoJf2
qReFUZ/Yoj1psMD8i/K3Mtr15q5fKkNq0AoGZ9ao1LDCC+56zQ5V1X/Za1HqMylDcHlYsfn7aPyz
NHR9sDd+81hm1Q61pnJfqBDVDjKttPwjzdYve6AgqkVjYbQQA5YFmwSrsZEnaPTmcYFuz6fxOEqY
qZfGuGLFiuVUCxIpmBuRIiDvrjeH7/RNVfEd2F74125K9GBOT4tF0gLgtVdXHxAg6M75tqmWYb9O
NkLFrqsn+ADi9lc7UxCoQ8zlIF+Id7vGWZcMezAV16TXI7B1l9Tm3pQaMnzTnKH2LUxpC2UHmq7c
ZvqZOXfJl5h1u76g0XZ/c4PTuMSnJZdpxOZacqS5JAab0F0lKWULWrxLjpT/5WPPR63X5q7o1xku
OHlFb0kz3LXml7l9XzcqWwD8kmv5sjhVznOd1uzGKhErW0xruNssTKA28ZKkok9Hg3YMJd24GU26
urwucM3kLvQGaBsyY1QeGFg7dZPd3tomnehFSwlG5EuU604M08sef7Rs/TS/4XlKzm305OlOx4xu
k6CDcwWLZT/9fWEtMtgnTjYWrr8cjN0Q87g5NqpdHpTpoxpe5S+ZhiutpaxcNfL/HE32uTBqMwVc
qgRdi6Yjrslx3b9+JS2I4iO9TiPNu20O4/4aQUExceoYGR79I2Zq+EY6DtnOE7+qpKSGY9atPE7d
LIqiInSTl5aOAl5WRSygENg0HibiVfdWX4ODKL8p5IXAXPc8NljFsUY957Z4WgBtEYryxhuIEy/b
OmiuZQy4OfK25ojtuHFK8zMOioth2jXW6PTNUqrKifcWUwRR5SMhrs3+WDFrO8aCy4uDTeAOZgts
Ut3je7qHnoRJ3G+1BbglVW0y4ok/iy6Ep3EyKQ/Sz0sye0Y8Bt2qeDR2P3rZc6kmpaQcpMOFDf7Q
zICN2kF0PqqhkqSVZchfqG7ej0Ze2gvI1rb8ULCsJ0Tqw5BUeLQL+hSIIFHZ8PbDVcFHVggQ3uOP
2i3wZuqvola3tjMQm1VEPLjYGGCZtfbloq2mquc8zciQMZMxTc8Y15cO9UT73tpqRYC8iS1ZzNdp
FaSPzt3IKVe6A6zodZmlZlCVCC8L14jZT/X94gq7zV4QgFbeO2oLV2XZjGxyNml6AnPR8uTgfx+0
P5NCTBFXadgPez/15yrQHukoAZcxc6Bm/gVywliqpMDlw3KL1raQ4hMQ9/+V70ji9RzF6YUEl35F
rI64mrE4eD3ujhYVLxRVycgFHDjfcSNVjxqrJ5kqCXPdvgPuEQnuPtohOcoJXMfpDblFq4oy0Pkc
bv2eqvbo6lKsDoZhMEdiKy5AeEtPoVYuZ0k55VAfny7w6twNksITsvn+GyF8KNzYE44kLrY/6vSi
wo3ZeNUsA8AiIKNxUc0O1XzYBMlO9gcjrazU96euM8g/mt4oNz/DAe1cbuCaHar4lqoL5ClDsBEh
Ne7Qcz+S48zs2NLLgyBZ6Iy/XEVXs15YXqQUf9hHJiuZh6QJBikUmUwlEEdrv9D7MRsN2BRPNAML
WR9rziRx4LwrI8prIP8sgvtkmh40XzXhS73XDFFa73pKaM2ynSBFXA2DKhpeykqQ+gWBvA3fyCCr
unSzB25VmrpTSpPKsgKfeu3KIQ/QCIDqssOhW8lHcdgXJtEFqWxkny9XKf34IPjVtzDYIBr6xeoY
qNhyF0V1UxLMnnPXfceWO9qDf6XvuZyDM+cofPKJekNv2tOXNsb/OeZwQ5210u8oVGFEOlq2o0MZ
BDMcPn13Xr4+MpEV+wB/Z7vAacua+dMOOdI85HpzBP/9vISs2FofxRBOqhr+haXFaZuqS4W5Ce5R
yAdv4G00iOhHkpkWcJU7Q+3ZvRzhzZkkcA1TR9V3+8eQNotI3TfnZWa9P74AnuV3qx8viN8pB5rb
QP1fonRCQrEftCpTAgRBASNXOcrH0FhJ7Ro6yDJ5Hpob1Peq+B9oVXEzaq0DPsrdSwUU7thwjjJO
7UoOF3WXEcQ9gL4NDZc6TC50QZHMmPHaUsW4jBac41+IBdwuxJSlc9EkCcndrBSNXAyD+a0pNpqE
i7apSgegyg23WWySDsLDtsXLsrIVFvk3SHN/gy6QtH06Mbs6VvIxtxHH5oS+ODIXUGBbKOYpqs/y
PO94S/+peFSUZlGjsnE2QkmUr7LsRUS+EA/jGwNDsOeGeFJN44KIB60/vGlh608SmphnMiWVlIjo
73eJgrAiRUZ5HnRAy8IGlIDdIAQeW+YrBgw/4RLFkikbRBzgwAtLVc/JVFZse2rPXH6MmNnEIPb0
A1zi3/kS+uhvffVP6EhvQhazM/crYqMKHceu3FHdACBckvT2b1c1B3mSvJln3Jsh6Pxa/jvJYTS1
b7sj+ZzX7u81X+Sx18Ha4GwUoRTBazFTIyNYTnnrVgVfY2Oak/p5zZJemaVLvN+7nNZkz2I09DCl
GzRzgANB1Tyf1U2stT9CRIYBBM68Z4xEDUAdw+os5xqMhcbNm0VZmcQUkvzeCknGNOiZ7gN+aEck
h0rBR9Ll5VCprcOqJSeW2dq+YXK82uWmr/pJ76GtY5PG91vJM3XEF17l6pWpCvIMyNXOzFgr0UmI
hCuPmSH8Sbdc7Wm4noiuWIx7akpOW3Yf5/9UjOP0hwy999ac3Oqf1Ji7+yMJdx6ZyiSRhBSSNs/N
rAHhIe9VmIM4bjnz3zEhe5TbuUSUDdxQV9n+6di0XH2OcD9vBE8FnxMhZxnQLf7DhFznlIU1Su5A
JdqHCcosezLelppyNcgj6FCBTxwDDyjeCJOBR5ra1Tt3pqqYcx7YM8JbB57NPcgK8OqjbR99Josa
sMVXTvTC5cUi7cy9XWu2hKcPEyuTRVakvdcZcEy5/BZksnsvz4RwFjwoobiUXzMJljHCxaoa8/h/
kGsdMnEC9Zs5LNS/X2AWy/vX0jRXvQFibfTRLdhAmSIM0fIyNd5iYGsWVYjbYvx+oqieucsaqcxY
nnsA+W9yyDH2SSWH/W/tQOOs4vJ64hipgRKa6MozvTMs6e3mXPvRP2aHGpI9VW2NsqWYMhrAZTuR
wV3qoXtf6GBPhhon8iqSYCa6uyUGDyWVaYhpN6tudqwNTNy5fsmZUAb83ye86bx9cbGQVkulrTDf
um1qXIuGTd71OyMhx2vaDni2CN2GmdeRA/08rxECTPsQzX+WK7nlXc7BFUEqCnqWgY7TMG63D26G
k5GDeGMLegTdcx+PP21pwOcuy0n3GcGkTE4byBBAtoYEx62e14DxuXBBtwA9LShQb8tTa0O2u0aE
WbscC2CUUL23HOp/vOzR+jpsf6KY5+Rl2cVa/PwHZLP5T8dabB//vzo1XV7nRnpK0uHHv/7Diml9
eZWvfkUdJ86KFQDt8o56AECpMIsnBqoDd33Nxh0o6CXfftDsNDlL84BZ7jbPRIZS5VGNy3lMethH
/pfwbTSD81qpkriYgBOElLJgLETFvjc2rUvc7iXaxow9i9we4CrCyxuW93m1wEmIjfWVyzLdRvVG
LGOoHCPqY137qmZETWUW7G3NW3xJI2p56aV7Ovj+KIC7xCHShUxZ9ht/cqS/RysZIhSvdRbOiDB5
cx7fvcuTYakQsIzO/0f9q6T4TvmvQzXV7WBt34SNxWX4hzhtWRNatKflWnGvp51OoBWiHzcC/u9F
1t+qLtP8rbeAz3Iuwc93RJwD+RoD3mImltZENmQeF9oP05WYhmddTFbgUqK9GadHJnvJsv9jxMdd
zPXPN7UwhT5QEC/bd3S+1FtvmoltcGVpMo8F/7j6ywIZ/2r2QxZ1c1ddOzeynPVBNdMK55z3S93P
8fcqzYcYGeJWYL1jNIFx4NpGDN4DXJPWin2849kL+c9MkEfxG8zPftgHvUpXpdJOHDgVvr1W1rzC
MtvJVv0I7xC1BchCvXKj7nB2NFs6w2aPbu+sQk1dvF/GGjY5ymKCgWBEFTYzij+xgUzU0ZU01twk
MJX5pwWB7Wq/3U3C3m/0UkC8TkLItXFXZkedJ+DYd7c1sIH6I0rgVogZleTrZj7Tnndi1OFgUbQx
MNo55WhuAH4IC0XmZCpAp0stTDKI6sxSGkAr5kuCrPzuhPWfK0wRIlwgwt1zk6k8T0ScTIGOh3+m
pF1/MHqDsbw6/f0RonHzw5IvzrLkPaSJSseEIFljp+PAA7afKX7pDzn/R0JF6q3VONUAubqIMEVs
tWgmlkzhh5KX10+NIG/iEhfSZraq5DEfCXr01K2iI3OYX0shC8GHOmZ537dkhiSrGzTK9hGg5Fs1
xS/gYFTw8dqqL2NCWoa843WxFHeXMmdyublPBS7G6YjpDJ5G5lRqRSo/qGZzvu6JEs7lw1X1280T
Eo1QpG5kP3tZbYgl4ReCyga+ND4CoYLgthIO7XznrhoHHrUG/NifX6Fso4DpUWYIzTuDd/vVgrCF
apsWTECnQLQVjdWy5plRp4s1ZkYhErioRzV1XKipWFRKHotTf98CHNdbLOnGeWxDdKlS7ZVQmgvy
AF/aYbHOl1YJhD9Rm/iYMYptTBgyCA3axXH/ZKKjtidBEYV2A1Ed+w0xZrh73mw64zy7jXF/gEEF
euD95SFz4cN3pwONRVwQ2shtgtwDgFrWVz9amZjEfWHHEWNM7vGbOMG/Mh+20Hw9zEIs+ve+y8XO
NiOWWx2sVjEswjv1GhXd7eFvJKV7/HGPH3Md+QhIEMf1dcj6ptQchQuUokcs9PsVvQkLgEjNdy77
nyhR7GjZxKm9wnmyiJTtrmXti093XsxXmRahjUwHzaEyBvcozcwfs4jvK5e+rG2xR+OYl1PQYA5G
4+9XWUrEwsn6OYr1zAjL5AMthCjfJj3xlAylliZGnN9brvw40caRcyVWjg1J79eXgAxLO6B30os7
qYYZsARrdmS6Qgg1L46tAXkdO4Oct2QXcYmJB5CZPIGMPjNQ0CWHnqAUUycqJASmMQjZKWVLnQSM
cT29GpayUBR6IDA0fO0myrGzs7qbUPfnGspczrKpB3ou76GmXFHJSA0k5uNyUu651mm2NwQlvSwx
T/g6eYcXW7lT7QgncdI6a3WzLcfvIHTp8+BfeLrBp6zqOX+KphfYy5U4H8dlexrG5VdUQGTvnjMk
wvBP5jnlpkKJwvJe+xNZwQyw5bF+w6wpc9CGRNiT6cErK76aBc/Uh7JHRS+R+G/wEhHnfiycBI5N
iw2GlfAbm0cGJ9ERSvYEQut6DDsO0fu4OgVZ/9OrAXKvsNcJJwRTMJ8bf8go14lM1h8B7k1+QI8S
FsIC4iPSx4Go7VBBqH2ebgKisPhavC24KKGmOM+C1OVHaYXSgjB+uU2NgXHhzI5OwDIgrF0W4SEM
FvnBVJOCLoEY7x0toRpLmEIFvjojlIQANTfWdV56neaw7tK07UDTLFdchb1YrF3TzGTaZeGtV2ks
VH7t+TGy/nL7RyLykMmqJCyEKMOZqCPJum9+nl0uqhKtNYRz179uL17S9JdWQ79dN1PczGPF7fqO
PMN3Tkw6HOkhUNnfasGkvsZa97rMuEPhaEFBSNkzfnhUD/rP1Ee5g/UkqnkamBXQ9gt+TqUR8u9p
hyUSwK4FwrnSFy1UNdY4dlyIgz007HuTiuubxArAzuc4fcdfvDFZRRl21MSOzs+8NnbSEHpm0LMN
jWTM0pPO5/T6XaJV+gUnq+EKU0W3E6nlnqC/Pv9vPSEbMR5+LH6aoaBhg1+OVrHTQ3XukRxBSmbv
aGG9n3t8IuGvdwJUVIyJNCiWImvZsT2S05VVUdfwoLNXmbfYo4Uul7wIRW9IGtaKLGxfear5hd5n
RBfekL8agweO9N17TlY7uQCPQ8/LJnQsC6RiXbuly8KNZWmXK58F09DxHnv3xj/BxTpQQjL/BaoV
a1xUMErnPMxT7akH+1K8DeVNxozkhkMHQ5yRa3aYXrK7ZtGUHwHqV6xzIJo8KRuzBkwFqLSCTTG/
C4uUxL9yK188XI/f7xVw6KAmWD5ukV8gC6uI0jQEZJKBUhS4GoORxj+8MipcGPwO5PziNAOatPG5
mRzEF2BHddkBNW2m+IMf9J29F7cF00oVTMUmgafQNrWNWLXeZbUdE8bSHHWW36+dNSweSXLnOqu8
UfeRqO2uG81L19gxORWYfTV65LXKkPUq7oLc5pB1EehRqwBMA6cC2gZ1RvAPHGT9ml3wqjqP5n7O
q7OMI7GFrMZCn19ihKVXuyJ8Wcejk3FtyfMKmCt9PKvxNBQvAfT07S+QIaObjhl6GI/csHY9nkGN
XExNN5s9oJuBOTvrFSE+h2/0HOCARVM8Rk5zd5WJcs47yvG9kWNPkyZEu70q024N5Beq0uwKGAnQ
3Up9W2/F9GiOXZ6kggy7gFntKcqIVQXnJLeN6iPMCU6vxs4Y4y2gLXnkJqaM66wPKEdR62Ais4Fu
3d+Ug2Q8VOAqH+j+fHoEFPBraDQgDC0OEp1QHesrNZTknMMP2rvDTnMADe0BEJFPbPYX3k/MVSYx
1QNhw81H5wEM+QRCS8iW+O8VX9Un2BxNx4jEFq3WzeMoIDm7JuowUQn6VE4XNp6ndTp8ylnoKJZY
VYVHQeG60c8MU4bNUZCTxEPvCP1Zf2ahob6QdVJF5rNU85kV7IXmZ40baJKAtix8ljD8CUhk1rKc
VHgMw0OGAwOW1q6mE1PMde484LnSDwKaKul7TRyAIzer5OIcvHHtqLDwwO58EPlrF7sWuf0GLKj5
Vjcud7OzvS4G7pXvtmUrx3ioY5tBABFGyFDFkUjoM1k78PLqBfZcTJCLg9NiEY1PF4KyuurIk5AC
ji5a2XGtBcF+KKtMHHxIcPFHCvC/FxrCnfIH5X8basgkX4Hi6aPFziA1G6USaSVpK5Iq3UJGLm8i
Sxidx2lCAD4AFogOrElbJFqtXSyo/M4IutU5dbxHUAskHApku9yE74u4cuDM5wthZSFui5g95Ipl
C4Khl4iI+c2zR2jCzb3tRus8nNJnNqyKVj70P4jAFVQWB4jPwJdrUImNif2j9WWnUIheU66c8/kk
I/FS3G9gUlDDM8u+JAwE5ys1uForfUGITfRONlWuqBy6kMiX3o2hmqF0AbIwF1sQ2Y95BJJmULS1
gt/3S5GPfaO2bPWdBy9tCDwVj9br71IzPjNylRJXC+s/+ibirJSNC6shVpW80P60k2sLFPMgxqQx
qK4eMYsTNOc0K9pwLCpL8MffOupJZOZhDmX5AtACmCBxD4FWJAzzeAZjKPftpaurRTb2G1e2VzGp
o+uEOYWoEeQ/9SsvEx9wqZG5y9Lips/DVHBTemnCj2Ws1Xhh/8QQOyBpJnALFmQAwTpEMa+TYzoQ
1DGs0RXcgRLlLk3k+m7etb/Ccpwis+APaJhqX7idXz0nLpKn31J14S+ep3ObYqoaN6sS9QK2Qvcg
hZ+driWor9o2RzrMPr15h/neFEppABfppQefxidRgHS4ETzCDOv53urRPYwDGCvkGtVpTtXgJSzA
N1yijueKWq2ob5fF/qEhraypLUDzm6nXVAdhN+JfIZmF+BbZ/0Grq/TlsmongRbsz+ONg6dJzXEP
NhodoyoYChpwCIdxDWg5MPmgnU5ZW1VRRtXlyLt0GeucO8QXAIjw9DGeqHxdhgoEPVDkMESt5zg7
APtcPIa99K92Rh9uVUB55Pqj5633of1uAVEUdC3k100KfZ9X9QG/55Zwu3qX7H+n2HyRk3GAyuhb
cSOFR22/7353hzfVrAY9CYj9Rd+okm4+YHca1tPKjccqb1DdUzImYrPUvbSShkzSSplS1i6wYSKX
FjlTTe4Mqm3roxxv6U2newlO3r16AJiqxIvhH+j0X4zgBbKGKHD6ZQuELemk9fKffesApnsZicWI
k+/gtiAfJ6Hc3aQsCkvneVu1AaruD9SWXu0vfocQZYlw01EUb2Z28D5Bme7YGPlKBiaEc5Do0E93
3O7JQT2fO2AbAYmeEmEqNaH8YFdLBsRYPKP9ewTzcr5ItJKD7GwLYae56GDXP2t/JiyyvnlTIyMo
XBpnK4m3Jjt+/AizNiPWzCqHn298sdZJDd2W0KGy4shYGavDPfBvgd3lrQgAQ9HCW9Tr+CuijW+N
hEGxfis5wk3jGM76yVaHDEnnkBS5wEmNumByvQGBwGaknpz/0WBDigpthqpVcJYSUv3GlMl2+q7V
Jl8r1oxzi84Zk7uzzNNkSxrVx3pWyIqQpyC3kGySDgEsOy22pYQ0ZU34UTZp3XNLMTXxu8PIrRio
DG0oXyn/P5tidFjnYV4un+cMnLjfsTG16SC19AUtfOh4SlKDsvbb9/2VeyG5HzvCyHvGuukFZCJq
780kdua6QQi3WoGr2af+5k5ZGXaBPvh/8SAdW/yGBGIOpNLsJ+IO6CTYz+2GRzP8SDLObL4hrZ76
2UawBfYeUzPLaaULwA8/HGdv5TwPB8NG489Pcd10c+KA5HsUOkFPVc548kdciAfqvzBJsMXtMq0t
6kgxuaI/DnPDNV/7Si8Yka+TmI/8u5u9KI/RFuo1u44efEWaC7pnvWpoLsIWL1zrqREKmA1qgXcr
8wOTfL8U8Au4btjGg1e83xco8bPjIXx9BY5H4QmsuZr2le2p3sZ0qimuEZIUzNgSLnxB5B46a9XO
qumrMz+fsHtijh6p3zrdHkms6QAr0Ta402B3YkFbszaejNRMeErt9idbFfSweV7DFTJtddALhAZC
Q4PpS3AcnS5Paz52F+ecOsk+pHcEr5697Xxb4PWR8JcARfl9ibj7VkW4esQRDWU0DUt0nw4Yqhu2
dO+8G0TG8FLymo90JVYmSKu3/9uBUZ2XxitW6k3me2jRrDSgorNMnBhIOlLLHOY26XCxYxOX0ZaO
JBPqpBREH+e1U+ZnjF1FA2naurL4DE135QMNKzBFBUSjEah5zDxBmY30dk9IrBtLd+z9IV2jRGzT
iMdbjz6Bi3lpgoQfaOrF2szYwuFiRY1dlmcnHfXoysg6lcedXJYp2OClvC9zUsoGR6FIUeijHR7X
mlh0P+Gy/+cFFT+9aphf1z0rilA4g3A+PZGnzD5RYGU0fgnwbx5Narw22Gf+PXswVTmmtFRC92y7
8F+VVdrfi5iW7yZcnjt11aYQ1j+h/yRG5EVnFT1MJFNMnExT6u1zvNrf+9aYZxDyAuCOsXbV2EOr
RcNpdRzYvY5T31pzw1A3FOHbayeY2iNAZVr0NzIEI8sZg9uNUqH+jR7utMPJh9RJCKM7fr6RQOhq
yTe9K9mhXYzOIv50Ulipn43BvDztap4dC+dsoZgC+O/Ad+fX1RuvEfLLrIOJbU8HSAKzbpnNaEw9
4lAoneEdXkLUIR+ZP54Wu7Prhs++W2JwfSjP4JLLg8EhJek/XbLntrU04wJjdj27gwCj966g0czG
M72820/2YHAvaqNthnDTt2UajlXy/G4V+ka4ds/DKcHuJDFfpx/V04YOGZENo4EKJao9gWLkv6U8
LmAfjYaWAPx5VSj9diSXBZ3/Cav351m9m+CVP4N5nLTgX5ath4Hq4Y3sSjnnIG/uG1Y1/r/qlhhv
S69F6Cfu0+1QcpwcTj6XcfIfi4VJXZZTYVn4s1+kNBQvKRuETg+zmkvdy1P8k0HChtmvaIwZWwq2
w38fa8ZS6yQ8HelZYIB77qo5rKp+JEiJTFXpNBp9qmh73gJoz6NOJR2PNU4USvf4yK60ER3wgayd
7hC0y6nKAppw9J9BqHqLtRw01Ks3jtTi8dpwmrh7iKJEy0PHlFkJQjaubmB9lAMdUuirWyHuI6zL
WcVEuMRWovXPFr4OplEIf8d2enpEMEIyHfF5bKhLvemwKnJmW7jgWm3JYV1QBHzTCkhDrv2QJsVp
cZi9TAk9+f9Yvi4iMx4vCbe+S/NRzApKHWm9EdMh4w/XqkDcwVucalEEFFOqVG9hsvGEUeemDCvb
cy6myeoZqR247o6if2dYlunfLUBkxiPHySoM+DPtPEOfM3UuVdhgdqh6KJccKC+Eh6PR3cJZm6Qi
+kfXaxmibl3fbCDokRPOJsmpZ86brr1d3qDxA3DH8T1M4epfwchDAt7wMCMJ8SonImPF4UNkd5w1
v4o9DYpcioZMF3zaHlYE4TcwyuSBMCBpTRhPBd/+J8KAyyfMCt/l+uD4+r4AvOQItV/rxGlFwr+w
qg9vrebJJVXLQq7pqWKfrK4RvDuRb08/gaWiCelibgvVJeqEXA4B7dttc3NmwtuDbjMk0/j4w5I8
CJMEgCdIAHgjhNvUnoySEMhU1goo+IXQ5tr4KJMLIdJUGleJwA/lnVYuGDL/HXHr221zXtEcM1A7
/t+pYWWNMW8gHXYxJIct7sV9s7wmoJBDUGzuJVNT5kcXbVCHygpjhI08D4rHQ/YbJMVbX2hqih6o
MEVsJIDs1XXaxNMCk5e5iScuvvoQEOdlKWfYByY++h6RRv81w+NmveX9Xi8h5U3EY6JmofT/44FT
Uvjs5kGPO47ovLh9SJ61pPtdMWxYpPXik+tbTXIdb2K83W0TPReckBb99l38lbA+iC2+hY16ZoSi
h3j71st9fjMCQtrJxBWbVIfzBKxwb5+RVq+R9J8u9xYorpNQE9Go0g2XIGhnGXn1nFlYY7/7U/sb
HxsdshNPOYpco28DgsCyK+L5oSBs4yb1HiUfIVPLlrZZIF+mB4yIIptkWezWZ3uOiAHDqCozBCUi
Sph2S5eV0cSKIVnG9AjPxiOS2MAoLphSuxrPP/lA13bQpxNQkDoHAVwHEoNkUsYMTxkRLuDlVsj7
/CrCNfwCx/oSr9Rr3raXMwYQHttRn/vLK3CDC9driC1O4S35vi1Ld2Ntw6Wa8cEjosudT9p7tk8D
BHbpfwdcUqnLYGDZ2UDX1ZtYZC45Sgzg4S1+aWCdy6W0wkfH21o2ZJzTxe9mvX/rvjhnTQrYd9E/
U62lpvx5lYn0RB1FQAFApGFh3v/KbYSud0ljhyxwkEVVJjMdIId0y+dbS//G1VNyCK10OEBBDk3D
HGednKyKOLROmckvikokyHnOojTHlGDq/qLdckcfnoH0yoSOQdx5mzpsNKmEF7FA4uM/cZD+5XIM
kAe4RtUASTijOA3z2kZqC8RKLAI+8ff/5AD/0CIJaX99DMVn3bQRjLxGbJMcSahVvUqJYQs7PygM
dLOXUs1oNPEiCZ7wVVCzpj0I1Cgp13ekeGYVMRbHLZGiKRckMQ2TqhP9go8jSkwmRGW27jNuavdt
Qan9SY0GRn2jQJS2wWZLT0IvmYY3d0+K4fEn6mM1y4sRrDbYSDCWmhXxiiksg9Kby15q2q3nIXGy
qPShtOdUVHKyHWYvGo6Ya9oj1HVedX86eemO9XeO7Fhgx+KJUvGyQtGm+I2+pZFZb74v/TEql9yd
/WChPbIbYXzcosDFfmKuedO1gFTd5z31GTfEaUWTH9N6b//dTaKDI7dZ/5ipJSY4piJR0UwtAqNE
1Y12S3m1+Io1iXHqdoDgHLUlJRsjVZgiy/RpnoqxfFiRkgvKceW+vRqozShrP1MRJUsXaONVWb/e
aLmELKHuPXm+c1tvMwhp7yn/mHURMzIiWWTvCy5KQAMOLSaKujnjXQvsbQDkensFJVnuCZogcsPR
1ikAWFs1pLcNy6JSDH7fxhmpl+hSStxn1m0QjqGr7B93z2JN3EKctGYgz5hUGy11R/LJ9d7Ppix2
iFZWG9mwAC2A1p0XEfyr50/KjwCem1ShuvwvJqHj4NHkq6b/wPMz3utpYsZxNiHuWArutKoqi96s
y5kB4uj72Cys89sL5cBaP4EB0NCfSVLNQL8DrGZzotZDFIXnNbfr6YqSmB8+GBopdANeTya8nKfd
qqFBIqoJltnoiDo7pTsnzT7zHi3WAIAZMwoHp10aIiJA1We/nYxlXorzUEMs4IVUsLZRpyaH+9J/
15U2FwsZpiVnNgtJzsCetsJsydB7O8sv3Fk1W/OmK7uVTwzGf9O2d7kkT8MGNy8JiJERKA/qgVLB
DkGTewiuLjUyIGHxbGhzjiBDGdi/Tu11pibYm/j2H00ClWWJqaYhpnfUcOFNUatdvPT0ZFqHV7Qr
v1+BKGg9/DwyXLiKgfAzvGTdKBj5t60ZTGyiCqPt2Gw9fq+Xbx/jO0Q3hxOMYG8N+KlG7r3sSF2a
E0Cdnted1xmkUIMRZPXSObFcBK+7Fm/M5zBQSPfusOKFAlY2q7DKhpSXHr24a00KpzpNWy4n+4ub
rDAYxEx88bpDjuHsduzT6V08AXDBFG/7dvWrZpLekiaw6it1910HopijvmReTlfDsEWtcUdbJgnE
u6AZdtwIIy7GP1jkLhzl4t9cQcxjSwe1nnTF8ojEU4nwMNZratisnNimdP5tJl/6CsS6AWuhTPgj
LInuj9pQybQadOMWK2Bi7uH5jkAFHLH7dVqmvjD9xFkRiIzI9bpyE+T+q9Hk7bSGlTSthwmplj9I
NUHsSxoI9pheizv0UCBD49zNZ42lXEqBSrQFAJPqiK210ZAoZENw6zZjFyk5PxhDgcVzt48UiT8Z
Ang04Gm81EL5GV2z82tE8BAryIxIMSzUP4o5754lBNK2V3pgUBC7UgRzPYIB/MEK+15Gm8HMMosj
j8bEm+e1VJk0T5+U6TazTVcKMS7kNMu+O1XAqvCSmCGt7NcKZGgU3bnel1TeI7irabAgldIGzPq8
9I4RNQy72eVp/xY1sFGkOsYjcwHgkU2CldvJfpK7+YqsyRhC6rrmVWLAKQVOqSqWMHaKB7Js4CI9
56j6Yg1eyPdE6tb7ULdIRY4feHCWsrwX4/W1O6yBZuxYA9Ban8fnxQUzJyGGJsL4QFFQKN5yEfcr
LElSocyEZ9HHHUE5ghnwytC9ZPWqMhKTkqqE9f2dZ6pgen80EMuW2GMaGOzILdQTzuzpGaCeVvNk
bIqb93C6ppKVlk135nNJXmiOft9+yOFtKU0L33qJwUmuhkRHeDUKQ7gLF0Z4K6QMRt644OuEM8Up
bSAqhP9WZvKbCtwb0kABllGr+A5JwAr5cQsrNQhBow+H4kmtjsJzxgY85WdC0+8lEKsVsUCQIHr9
gV8PSn/NdLUm75MxtLG4kXR6bjYpCuwKFJsB92xugvzAUSokgzdc8WH7R96nbpowvTl8IPHVbxjv
Y2xWIL+ovfggfc6UzjNa+E/aUDGknBPRTCDsKqL/v5IGnHtmkCaPzSx+mrjazxBhkes0auJBvGGX
PMVi/SBCBvP8ew29DRzXSEUDSLWrYYgfm3EFciHuNlFFDtnl5CnpcqSfkHdNnRHvXBdIIAmVwLD0
11/7CHPBv8PKmH3GQLBx9MA96IWateYP+Hk353+ItLulZ5b8eUG588z3RDORtiOa+KyW8UNJgwj2
BnNYC3JWQW3ubUamvLGJ0A8Xt9mzjhvt/qWddRQhNDBv6NQpL4+P8u4gfsuapNGVXlEKdnga0BbQ
2d3jkMMZA1NcubgGGA0GQ2hcC69Sp9YUelrlEwFlfKU+gzqhc8hypae25RgFlfnjhwi4oRVdRDgm
M02uydZISIyuNEzuNtVoVOd+XGrLW8GKZFsEnbcNcsquBdgIHrftKiPjC46YisjnLPecTksz0h5E
pzdSLen2M0zvb+AUM4yLZCcevTvK/lA8csmytvqSH4ykU2gToGHOW34SmLOgT+kTLfAcUIo6jJCF
R3qTPsDThwGOUe2yMmv/q+gFheZNaRbzeD32jfuCl+0qCWfl9UJotfhsAXsOLuXMQV1wf13lATam
HKZgoLutuliCi1nalefTuksNyY+PsABIHkcdX0I6vOsDdwJIb5V8L+QD+MY86nW2jT2BkktgMp1M
9RRW9mCTGaeditnVNXaU3I6rS5VXAba5x9aC9wz0/AdSftNi/Cri2NbfOJZ4ivZfYYXPwQAJyc9P
ltYW2rmOxZGrju/9H4ne/oFG9WHW3B4OUvq/2svOEjElw4iO2dlR4cG9D7S9A1U9lN0fTLwHPuKZ
ijVHPCoICCWTxTtEClNnTFEl62RNzBiZNEqZjUENUk27QxDnuBNv+2pcHjKFSqjNipwWLQAiK29H
lw3Ux0fzauKrG8WvkwMGQmGHAqit3L+p5WRIU0zHQfXgDFqbmw+GOG1xdt7yEIhh776CapA9rCGD
PH/+FpgHJ4obCrSj0JeFAY3My9Vcrcc/7xRJ9XEh4Fky+jYZUvg5VAmwOrLjJ33xNfKlxEyEtBIc
w7IU/D3FSU3fAW1jBYVWQIMMiL1NLYyE4vvQyOUSnR90BFPHFhdd8YHCpa6bW9kJUaCgesr23bNk
W7P//wOD6SlTV53A+gi3q+lZ1s9/3S8bW8Ujc24g7KQ2khi/KLxJcJw1ZbSKMwmNDj1AOF/j3/pC
0l1aJgCpNqe5rrNncDvNqMR4vOJtf64j7J+Fhfmahvz+64Ht77kpVMDmYabsUcRcKpq3KWa0zZak
4cIU2blgW7/WZQVicpRFVI2/iC5s4s54OArHcTcav75Gq7owya1Q8sAQTZMCSVvcdUaQwjDNItD+
cfo++IRt769d9YhAlsuWbIg2FwhlwaNrOqDlyYSZscfO/xA5aSiPg4mQWQczLZsXhf261OfaNYn4
FaZSE2kzjLIsqJcXnOrSniB3IzVAI6xq7ua0nlYC91CfEp9w2VRqLsBvrwp2pmOa7WUpwpldWh0H
Oho/V43hVq/hDttZ9roHQtwSr58SO7JOJCxtjhMuZBv1d9t+SUq7Qgr4pdIY7smaiOSK6puKfCto
yFU2Qqjx23C+6cjQJySdVYZNK7/meQ9sZYnWNCfWHc4FtroQfxzhrvxCJ+AQBTe17NWqgxDYUXXh
mveaLFjC1+5hhafuomAcwOOJlVodfr7BgylDX+1h0S3HvtxbmnzBiGl7xzaTYw4Kop93eWeUMbdN
UvgTDkHJwPtQNh324JJatjUCEfslyQuV1p7PRZiTUI6dbxtobSASbnE1XZAPueYJCKB/s5h9LE1+
H3i0CQ4frN2a3qi8lbxg60XQo2n32iDMwjFS0GkfzvQKy/FXF3TfFtYJTufLxWOUwOgwo2bg7+CG
23e1QotuCw7a+eQkGicugXZ9DfaUKtRDRzR0O7htGcrh96EYkEHDvu7hVyFHpS8VGjxbxzhAYmKC
nk4RuWREP8E2hT4JmlMfE6S1PZ8d3YrwiMafYM3l8W39bxllfCXeTWtbNd6XwWuPSLrVys2H3coe
4ymrF0lH4XsVbDyqTgS4ohI+dOsfS7lT+8BBcb2jZTGfhpSepGn0kvhuYx7X8PrMAkn+44x+zMSk
Jn2tyVXEY/RpSTL6suzpKSTwJRJ+bKsmR29N4PQaoSORsxtZAbA8auAL2yl6WCF0B8xk9/glr65U
T+gKlIOfiDqbKwmyb+6gO/9hoX8i6TilXKEiJdqkBQGunb0sfOxh4Ery5C5UWgzFUAOVgos389o8
Lpzo2+MEQ22HeXxQVw3Vr+YPfxGiznwm3FM7HOwZgmcsm2MsqzAQBtaNgK8kvqmJPjISu/6WcDPL
KqpsQ0iNFB1BU96ZDmxYocGeCPpHgjtq9vcjSy/g6bfQcOq2u18m3hQE6A6o6Hmkj6h+rhr/KG4C
Rl55jgwi0BeHmFvJMcLCWUjZC9qoouP9+G668uhnZPmp1LISfYoESIClRTbaDgaS7uvoXzJuBBQD
kaEQhaLI0AaFa8WDXe/VUr24QPSBbWHfbKJA+4r9psIqlbeAzBalcS2K/BXrl6Jteu1vwrXRqdEK
8NxLj7iLlvkaFwWX8FYNsBWTBhCIMeF9PcUi4uHzFeOhSPQs9FviK2330qvATquqPCEsBV4pHbCg
ztOiK0R+MTifOi0iIKhUWYLzEl+ARRaWxY4WYQhIo9AtjjewKr0jjMyczLtUNLoRo5p32G3OuDK/
gD6T826yIqM4tw4JIVhraJLjW3/C+217KFWbGGbZizNkXv8ukRmfw7uOw/3XsdnRx1fdDDty5sbv
KmKgQm8NGYuOLb+zm5dkPnMkOOhTaI9++A3EA7FDo3/4v4RG7grBZu99JGuWuJjWrLbvE4GP0KdX
i5No073Fs1Cq4f885N9KMPN2seLY29X+totsBKMGrwJ02J+fk5lWcDtS8BlTB2u7VQfKBVfnCuHD
wWY+afqJd7WIqzWWHCWzN+RF5tmJnaOAhHeynm3c4umvKlRO7SLsoy/0L8xKIhgrS5InlqAjXFgv
IxCrli5MvNxGXjAb/OG/rflrIk//Sm/wLCnq41XMIqiLMJx0H6RbCxbJ1H5/KFLjeiT55Crx9wNT
1QwgFWLmEfKP6rlklzo+r90mhxj/7s00S5VXycLbWqYk4Ss2V8yrX7motYIN+DcHz5HUEByrUe79
khHz3W47Ls/uo7baSxWRpu/+y4JtvtLqRZoTnQtrk46H+xqMwdh7BzfAtjxSwMUCAOZpeBFv+3/Q
lP40OTXvjsZq+gsUi3eiszWd/6SLWgo0eTF0IakaUSdL1LOlMxiakcjetmUmM/WE74qq3E41ImrV
zadqDBDWm46joAGUpsffqf+NLnDm6NI8BQMyhT6bWd4fPiOjmMLfW7DtCUMzoclzRvn3cj82fN7c
odtptVm/IlED/7ThZ9jwQGYScGqDOQ3nP7Fv6+/gtSHNgk7+aHR/Vi3kIhF+Aqk8JIrT210lAXRm
Ay17pQYXlTCAqA7FTSBWW/4gW2MVT4DAZDfEhhPMhnqXummoD4TI12RXxw61u2Bu10kzSrCKF9z1
HShf4o3aOGuz4h3Nr/aE854H3lXc6cW2wvQSNcTSLRX9WZq2O442QPiZrT36xQvaNoZWdynHa6QV
3aFD3LirWiIWFFbDqKPnGPsD+ieCa+kllra9uNJEeQC4DgoGqfBs5s61s/vdiFoQH6nm+8wktlP0
age47R7yKtqce+BHeFiIuEHHp7HwuTSH666s+6jcassi6McMK6W1ByYV1fvMtlEZTnEdJwt9oeaz
9/Q8z7TMDSrHbCVGqxhhMPjpEzniSikq8zpA8UWnVRYcUmJFGP4J3hoDpTBIksPffMRmLjwdKDDl
I0hK8EAXZ16P7t10BaRPk6/dj4G+oPJVshYWY2I150ZtbOIaGAUjHG46XxMNnHvCfrBY0QHx7vZW
bEkglwxDo1MYLw2gYrOLpBshPsWlvTjnxjgluQxIOiOrWXmVM2iXpD17S4YhqrP85YWo7k35ofrp
4Ap8h8Iy/+gdEkjmHMA49I71RPJWFXWLmyZah5nBev/V0RcIWuXjshtfqmeeWZtEnrDTwWxTneqX
LEEbn+occJtJmreoQcS85FsqLz6Xr/6TD+Uo1JJ80ej+mTLW7wagoiKd6tGADBFKV31dO8oyVo9a
0WAD+P4HrdrVrvj5pfgNDCFuCH38GCiiP6q2p0ubtUyXeTm8uo1QklaBEL6SBVVDg7rIjVjKW3yt
499RCWmgCUFKgW382tfQ914OP709JaDJjUfvCLErySWCvIIoCnNSYoKOvv1UrsUK5NP/d2Av773W
ZXnY2fiKMZH7PFIna2IETvou2kcxVgnqoOrHas0cpiEmGqnFGeNCdT0trtWxu9goaTfRWy0b5LVk
XXlKzIjq5HUHYKfRvjodVR6ABqo/JewC1ac3zzhIZ30W/cTqaE1s+xMp4baAuzF0lLQdTlvWfy0+
DwS+vrHQWnXZhFjKzsfZhC2mr2TNfAczv7T2i8gLxXkAlTzcsR0GAAm42wG7mzh9UJKgXv+DlzHF
tpEiJqT2FCcmUU10keK38z8xvTv5Z+NeeS3skxfgwE1Mt/xtG68GIOsZYd+rE/TL75qgiAF4efw1
/qi4i5Mf+66T/eCoqQte7X29RUlDcxA9i77Q41dVdG/wPOHuc/cmgwfQXkpi8y7JHYb5QroQ1Z+T
+auU9v8RiHp5Aqffkg8ls6JgsoWsc9AwaqRl4dMqPgjC7geLVqX5j8p9KAFaTiRXb6wKr/X2YA5d
Io+CUrmqOd8BRx0uETrK6gls6J1RCaGSMtibTtvAKr/x7Io+8IZ1kyGlrE56OaLjtmrZr+3DooMF
8YxRinEJs/Z55x5zA73mX6PHG+m+O3DyqOt+Bzasfw316vMXbOCfmsH/jhBJ11Z0RVGoldziZQ87
sg1QQPlVR/zKaqLfM8vHNXBJNFH2crTROGbEsT9R43diNAeESBhKclT+xVSHrs06Pz20k8ulMZaO
+B2C1Djw3KOoOuUm334O2PG4eO2SYv5nBWjghRvmP3kORQn7W1VZM65hSgNRMbnKWvwFpV8xA2Nm
kZmqmI3dyt33p+1K8OBDqJiQ4FnOlPQfEajOgwjb7ECdparSVK4AKIrvh1WbgWxJZLz/KyGCXXun
PFelS1P649yGyL2opoiw8H6oVV4WYZV6DXOr/Z8rHMYVyz3AFace4njXg7AY3HE+47LgaeP4YgY1
Ag3Aj/CccbSeSNIuffAcW6LDKxZbWaYSg75nR9VBvc41ySjtscOnatZAtijL+aMyOjj2zMxrcKDz
lDZUGprKQFMtqyYhDXZM+IyIIpSSD9CnQojXfLMd+noC9CWpkUvMXJcXPqqtGE0CpjXDMkGluxZS
08iPunjF3ieyimaCMuR6sCSa+8BHFvvlwN6oOH1wGBoKJdk/q3LrU6r9g2vvlauCcXcpffXwqmTb
N3DTcpLT9Rnt0JV/rxZLkDL5sOy1xPzn0KJukObgMYgEP8Bj8IRqyGSyy38WjJGbqfmgrpEJxBZA
0Ij8u8d1BjBe8KIBCMT6eZZqYRHO4ix1JAfpGwERfAslvtH219Gc9Oy2cAzBaQz7q3OSbVrwVLld
L3TDJx7rKeyC6yDg1ZsG/N74BwJ6swjtHaBnCTMjKUXQiK+Gc8gG4a4GCDDZM4y4K3MWvu1Bh9Bo
IFsQru+8cq7+bkZ8301j5bMSbr1oHE6U1qspMTAGL2cmvXrR+JNFKHrIxBQ6i0z6ytMC5Y9DCQvd
wUYyJzPqkLCevMcf5jrYCURnFkg8y4FnVAQEG12Zmx91tKiObrODEOCB61jQ84HUTVISbUMTf5Qr
PGjlVDHsbQzYq+kx5WlKfKRjhmqPUb1ydwpIt9IYwPfU3PSmfqWB6TT9NM2keA1IbxgN44eVKwX5
zuTZEvJOF8i7vMWbmxoJbELl9vOmUGJ3QwNuLNFFcjyQFzEQmKjtHocaDHIOPuz90qd+fx77jH6E
axU2Dv37zb/PbI8lJFVMAfATeA6uEvqDPdAhgcnsCEo6NH0l+c4Vh2RdMCJEyjxi62l6okSqOCQh
amr6XP5GUHLz8xyiBV2k+w+sVf+Z6RXek7Fh2BKNhZBkMRzyhEHqQn6leqBiQYH2mN+b6CnbKgYQ
KK+mZXjGa4347WDe/fWZTtdGn+pQPRj67Mfksz2O0OANtuprfmoExCjQDjvUId+frEAKJ6kJUb5n
q8mZBXIEows5RV/x8h165/AQqF1IhIkwV05d+yRzZPVR4A7gVcaCNHK1rJoDbdVPdj0NprSLaAvU
LI0SM5q+f7hp3CBtbUU5WOtw8h4qacvCkYZ/Z+KKwQcnnV2yDw/OETL2Zs151f1AJG3fP/CLHbpr
euNGb5KB5901Lbtiq0JQbaIlRygN9qw2p5j8hLvBGS9RebEa1REANPB6IXZt21DIA0+IJmEkLROh
aH+DgtUZN+F3o82F8LP6DELJilX17vQeQNgbxZWSJiPxYUeGarDqAul/nhNeL2rHefED2jq4boav
/oyqlhjsw1QOcj2/zPqR1SoMlLmgglIWm+9U0P4Bg3O2J0bhQjb+/UYWD/qKtE7zviNp3ryx76xo
n1+j8f+Olk+a3L8pvdTVy2XyfNAjloi3VFtxUuQN5vbXQazv0w/VOIE501dZfOpUaOiagx1zPrb5
nnSjXAvmU5bXTKpr9Xut3H0/F/oTQ+bbNW19xCPHjDBssvlbSTfkeEn3VrLKvrLrUJ6cYxRYRv/v
wfrxf7Tdtfw9vWrZH+M4/oAlHdgYkgWkh73IJku/MOcESmly/WxY9L0lKu3Tzt7MJ/ju9v7ZV3k9
P1i9q8YNdhRpaSOw7qKq0WEmeAlVRmkRiJHZ9XAdQIYy5g59MZOa7QppkRBx0wvewgRkmSGwN9JM
R6uhXXfMk10jrPQaDiSY7qI0wO1bq1FUmTuoaI+aseEitGS5rjVNc9mlibZuRUahmOclwNYs+59D
lT5wh21w06vOcqf3pE+Xux2/2rI2B7h/9gZEEYyWPNPy3d6wij5ol8iTJIuch6olZgBMI9bxUg7X
1d+ZK2sFh9dYhWC7w8r4yIAOZe4JxVz61pdj6NCVPM4xHZ9I0c4Xo3rAPZHpfTgpU18FSwtB5Eoz
DBRTlE5pri0tYM6I2aM8W/NXgwviHwg2gqGCdAYqvszG3pcv0o6sYNNxBH/aIRjWOzqvVuwoWubo
KJqXsDhj+HGqakDoVC56CR44/Qirj6qUm5QaWs/SS7OYUgv0NDfisOZVNMdsqiQCEdtHLkKy0lU8
K/xAZ11YZFKHF5BjNWpa+5wFUMPumb0dP0xEayAPR4iBdVrL+cBr8/5hdmvLnd0nM8FhaqyNGhwI
xfTiJA/bk0aaPQCXzyoZehUotR0E2N5yja/hXguS+GddCmqX6uwfBt25TERqfaJ6GJs3qgjEiAOU
O2JCcXa1ixjIVmMXOZppL57hNjsoAY6C9qlw0/zIzGQmv76a++4kDaEHYb462dKgxEbGM/q5+gbl
OdiZpPCSmGfRsvYy4eNKEuqpnH8Z4l7Cc9emruUH94ZTJiItt7FzABeeknqTxEM3a3wY6Xwl/fF8
cMd/PvE4axZ5Dy/E+4M6f56DMZygiYN+ON3hT9Cd3Z5PqwsDrvZ2h9g+5517MAOj2RpIkFOvW8Ej
tFHVhDfTiT2BKOL2vkjYPn1QVgNK636SKs5drDm/qMkdUDtE0qu2qbnoCJobi9I65zPqyYXgNq7X
A812GFkASFFxgRY7MNJS/7JRITPoqvGi/t9eeYS93ABvgamkw31J47IXi/1a+ZUhPRRMqsfDlBZI
9dea2FHjPDQ7160G4l81Be4BPja7u5nmeRDJGbG17jWBHxXe6zqCT4wCnP/maYO4zdDRMNcahh14
MCgeZR1uK96/dUuAsI5ObzKRiudYAAjizTBQdoyd21OXIHXhgTMwN1gpS2wDRJWlpcAB5D+4M3cQ
7kqbD/YnR0Y8FNsE7GaXYitSaLkgbXvU+mwqEiDnMflhZ16ijnCpcvDRJ9oZ+AjhIe/v6dpypuWy
FMnfKyxoyc+DinvhB5bHhPQpmXVfye1j5r4oHc7bxXKvis1uPx/utPSlK34bv4ZGmQ/YmGjPUIOw
gzhVQZpIkpSEdlKWo+vg4W2AzE5NoS93iLBjUItX79YP82xQU08MWINK/NVvy1eEiOPKNQWyHBKD
VZeH0hiZ9EqHrzz9joFFqfrw99c873aso0X8Xy655aE/z4r+V5RaGkck7VEbWwfJxnTBlWkvqNuD
Smdy0a4thlabnUV9ZudOz0r4+rZO18RO3UsVls1aMVyUq7xYPH3T21qWewLr5KqFoe7UnsgPTqYg
W/ZdxqmnCM0RPcHuNPalTjQKRS25PgTkZfxBf9x/NF5TBUScjL8qGSVo1rVjt4EQ/SCSXxzg6auE
ddIOMkABOYBKYmj/DT9vvfMup4aYUV4PVxoppaTtnZm4D1Ga/Rzsef6dPJrMpZMZGGpgruTXXwEg
y3o1r21/VZPi6iMsna+yK2o39WGmHu21Hos/jjRRSu+kvl1VgkExjvoHw6vF+jFRE/rfNMtMx+sV
E1pu6bcz2HI9Kw28QPay9cFnQu2m1CqJkXjWs6KFMaFjAWelJVLJKwl75t10Qby47Tc8gGb7XD/Y
dR2Dvgq6UCkp+KGZEiwgyiA5eM70K7i09bEuFPogdz4O8NYIm7YAlAcNLAWt6iTzHWymW379wbJx
PJku7dFgc4YpeG5SKFEGnmYqpkZeBuYCjPTDp4omShcxKECRlHU1gC4Y45eFo1ZcFbtHaCzXcW2Y
wUFtsnOxt9jrMTmypvl01W4Oi3FYhwb/HHwSBCDYdoCz1NEUt/ruOFwO+M6ioPlkSF0db2FMk+X9
OgmUk4Ne8rRGiJrFfckZ+v/LoxEh55xlX8B11qP/TFjFEgjH8LZmimn/VacDN+p4e35Bes7yBFQ8
7B34WZMKLxFHXkYshn1L8GWHHZXv0QrHEUsvq715Yy9jnl2OczIdHApvLKLrbaE/qJ0kj0VPJ7cF
vRBCFuRm4Wk64cnU4MKWQzX4g5iVSWky/I8kNWrO1Md6hK7DMK+BP83qI15PsUz0a1XGlsCdJHhR
4BvSDYtUQMm8kKvrbxyyN3HUOU9jvv2igRwgWGwYHXTnSipMqHTysUNM0C5wwkMFMcvtnfkf7flv
vdJXRSuPi8he0LlRAmnfZxNz6/yuwlHCFCwLUBAUOjJzM1ZO601tj7jipNQMwYEpk5uQCXJgSUOs
R28rM1VtBTX0jspgwog9HPjdTZVFvz/FvIB3bsHH3QPVZT+5jewyrEWC73DLhAKs46hjmWCop9Oo
TKESbyHkmUg9c0VAURBrzdaJcSiDIGd3Gvw14KWc6jegjPLU/w6AQ4tdCMsGo9tLIOL6Qahoo/ct
cppV+uazNh+wvVaDtvsK2JfnQ1bRM5ZsZKVRuEZwJxG0Sbf4pjwnmBKOboCT1hWOPGnRhbGiuz53
57FSisrOHsuSyxivT/a6BX2W4KUpCh8MY5sa1GjQKfet+8QHpOtfrY6VMgxrshnO6nHjD9KAQPbs
jdpqr5c9kVMLunHcx5jW0yn0iFl3/mR8K7qjStyaPxbPgrMikm66JH91DUGbUQwak0u8iUWTNhXJ
ujTsIAAVIt20UzP4OAHy+G9XQXhnYZFDtQBn6/zGV1GWzxI+0wEgkAk7TJuV8JpEQVKNdlkkbpuZ
awxFRuQBKJgOgCF8Mpoj47AutfWxZcwjCnt9dGgtMmPlEOiUeTtt7N+mzzVsGNA1WoaPNI7SmpcY
ZZ9GZ+qyN6IRSw/HLfkwxZIepkd1AqcEwYfg8y2ySibtylAp6HDMdiRFA56g8LYU70qtUuNmeUSU
l/1guhjt2CKV65NSczgT6z+Nk3S3WuVdRjYfwQVrjNywzZhy4ucZ7mBNbiKjMdTSbUemFNkgJqPj
3tIZYv+r5VpsUJ2JVNK8laOTYhjMguymuTJ3+yCSJd/D8TorS3bEhYGJ+J8MTPulTFifvUBY9cV3
IT21glhEsyJ4586LLImmXF+pM5c4xgzIWFbkGkvcXxnNXo7oDzCVl1HeMtMXh5xFXTJTl/gQiGxZ
NI88OntbcP92tn205DAxNGJA+mX7g3fBf4sfnHZXuKuLxRR/T1b1Rh8qV6axyiCROJKBZ355TgDp
s+B7MU2T1NmvVVLAceBsQZoRvgJ+l++8W1KNU6KTcWuflr6zgcJkW1vtopoAjTDXJ0jZxZ1kLU8S
gMCY5mE+M1zDFtec/89rg6XzMazhRk+7Zt3Ii5EC6ouNv/RLbu9nUqPpY/Ahf9qppw8XVsKGli7p
HEm4z2rPrYJW7RgDM6+AFdtl789ED+HPrgJ6l+i8eVdk4kw3Jph2oinXINtlMNWB6++pPthmKfHS
75QImlUdKPgQwre1Pkh9GRYpFZne8LcPfMAiiEzG22HF3fEwWzwWeCIyqGn3RGfpUVbywZPQgWtk
KohzhaEGxJN92bxi+0G9UEp10bXcKhbpsqHsKMfSumuyYDw/YDMMwxQnjsjM8XEqBan/qzkZ3Jfn
jIjNOe8oVf5SbuuWz240jSdEEkvzvrD/vaQsZDBat5OWD+BlBrz2D6RKMW8Zjw8J4JZoIp35n6k+
d5hA2Sz0vaYJp1960X+7OkI3/A1lzy+ZMkTP7AZyukAAwvWfr6U31zVg1tVT4QRlmwn1tX9UiYUR
wdPTgNniMcr7E14v4TB85hoHnebaWkOVCxQhuGCbQE6ukj2Fs2hbpRlfqZl/XMeO0FPQzaGpOYne
CCxKuuyjXX1VbgaixM+D2aYBfSz/paJaNCiSYQIabjuu7de6P8NxmS5qRx1VlUtZEmaUtA2Vmbau
ve3hd+KkTxF5Esh90SIzcvahMDDJcgrw0q0d8RBsqwte/0MS5usn5g4uqV3ISbCT+2z4R4a9KtYH
5qSghJZGApM99UMPoGS82H1R15jM83EOLuT66SJG9wwEIla8xoNGCYSmGlIffgh3fqy6kTcHpxsx
2wEiNTp5zTm89OpZXr3tWzm6jl3DjhRJNA3MwijrfwzqCQzNoevliA7LvkA3plD/nx2QXDISvfPn
CwiztFCHuZ97hkU6wdQRNlZe2MHhkYcu7sR0xF5mLdwGwRvsfZErBF+ZJRSQBpmMlrR5y4ww2C9H
kzgjQ6UhZfcesoEhVAqeN9q1AZ4QrZ7CN09LgifuyJx53TZTpxnSsKvpaV9NUYP2qhQtrb04Nwde
sUfnlXFqqquXx40p4/Rm426FNak3xNTIP03u7FiPZ4ZIIHPFV5lhJWpqYjoDIjW/mhwBA8X/lIEr
LYQui78M9wY+VaO0PxSBJ4IX7zfkLMOO8PEd6H7fyYROQGjbeUbKGGNaJK/0elKeqZIYyD6TUB9M
mhvCqd2QnAZTVpFbQpLVep47YNOKQYpjKe5HoPDS5xYi1E62nQO1qjiYa1cKhzGiAlE6mWI/P7DF
2+hZFyEos00DRmCQAEYYBIh4mEhabrBHW00zvlmVy0hbIXZei6JGXIrfLrQnkrJtOATA0b2E2010
DpZe4vL+nlWn/01q8KG3PEAwGUxKZBwN3FdPm6LpMrhep0qTmnf7dBXjrVhMBWiwgmMhzzpMsgKb
Y94G7Y3pjShebh2t+v3nwAijoDhvxM/j/BEMy1EjaburvXw//A1bDJHRQxnYNPkDQrJ3KM8HwpOI
bJ/lV2tq9RNQk6f3QFfNZlO1dwovwsqJeUVcOPceWTZUg2/ha+HefCHPxZMYdFlN4WoZ9hNj92ra
OsthVMUUC3Mcl5uIa5dGkd6TluVYirIbp2LufPUB4Ie2dSO3UxUBZeNCyN0UlDElIA9wqevQBvCM
+M039Z8dyiF4yL1YROn1AnBTyZbG1JfRAj64VmHfiBCJoWLPQ3TUIRk3+jha/fnNok0o/1eg/nB3
c+G6NJ/d4JVitehhEAdJJ3a7SUhSrReXTtFYvv1jzJGGd9TYwBvV8oYr2oIxT6PMsHXJE/rup+Id
3r06D5Zmk92FQBQGSOCL7Y6JBVYHiiMXdr2JZXRlzfNw+PKRYZdWE8eqvGWET6kdS7gIo/IESFL8
scjuZLmCYnCYF7Aj6cYhs+REQ0A5bmgVKF4hpEwrSlEoozxwqXFqsBX2bBzbjnpLSMPBCciRYxDx
6eBciajF78658WyyLmSoYBtOahK9agIenydZrTewj9cDlKos+bY8PMzNi8FlniwwHysPuaPUDy6I
wjsSxd7IqWyLCJH3S7n4UHyBS6u3cMaIQo02EUBeepmLCdTik4/tNsaiC352YJxGPYZqrT+SQ1Xh
JXMNKAyVfHgcFNKqKvc6+ml+cCyON6MIUXO4K2s1UOfHbWYK8QUCcyUVV+xorAInLqROOcZTQVEI
ouwDJru0gG/qQBZujcl56vM+d6Gg0fjGll2REW8yTSMKA8xB1A+i8FQTc27giC8iqhfnchQGiAEP
XopP4ZB/krO3BXcQnNJ+Vsia1okjQ5PxvROE+HD8IrllS/fxL0ymmvyexju3zqGGorls22ZKgaBz
dJBB+oTbGNWoIIAN0LJAJacAi3hVzA9aImCMTJST0cp05UwxE58J+8SvkQS+OjjaoV5eAIIppqds
kEvS09rvQi9dgZql2kN0AJ8n6eFt1ez5CyHoL8BBoOcw6LoPcvFc+LoRinYcpOUCN8u3aO27zaqW
0NSs8+sL4xsIQIZssO7bfuBi3xgc68vp9cvGXScl96YeabBdcs0NcWVqyMRotopCSWw/T0bBsXv9
3mQE+aQNFnYBmvCuk+NEeNbezGjnZaFLQI+lPlTXZFj7OafNuflYs8A0k2svah1jT+go3DWd9tx6
+s5ezSc4dSirkfNuJX62hV70YYQU+CfNSKolY3+uocJafDbcTSLFscSho9wqzHdO4gi1484F+VFD
gdO99yobDKVzrPcP19YoSP3PMBtZ4cPQTaq4O4Szxr4sQGnrLAtUJZHCZEjaD4OGtog0noQrYL9/
bAz15Db0pYA4AndEW7HKs1MMkXqU7tjA2yp9T9/KBW2wtaHtUF+nsKWp/mZ7KfqJVIAhgpKN5BS0
GolkEr9Gnb9lvijGSG9YQlF2BcCdZp8Udo68gxzp25/QchXCVa/gwRLckf2offcLrLtJzpPpFzHr
ksh2t0q+brfbvKNBg+jpB/oX9X7Y6gMjZ4RXdhsxEMn+7L5radZPmZZ5TkmYPJJf74z1VcbPHX5k
+NP5w7fQFD/bUXtH9Wtwk4KIaG8kSmikIOdtdatiGD8U5O5zEChL4/8VNFfQkuuzpEAdTtvkbcq0
TZLoCIwXoKNRDmmQ7j8rj0c9mo8JboYqqwr8Mobwf93sKgp216SWaYv6uj0MWdKXZWvUvJ0XkECb
Mr8QzXBO8TU7cDbOimcXY1Awi1yQB1J0ZhDR4BSM3RuU6jNb4NcbYdcWbYeHXCabXFBL6Mzz3RcB
QnbECbMh5446Ik0qIaYKd3IevyhztJLO2uKH4CkfevelX4BPYN9abfV5rytQxVYDFz3S5MAGkyoo
G0bFfUtEEWoBZ5biueIsAoZIXadJIjrEJQyE5lgCH/E6MbEOKo+E5rQxuoRoe/EqrqvWy1BGMQiB
LY1hKHZ8+hzz8xS1PhYV/8difL4gwHxLwOmg6S4JVJXAZmySngPpF+tzHtBNsWp9iFwh3wSeyUmt
JhJQp/UNCMWl415PSYCbl/TeabRNepW2xH0H9gq5UyAo6EA9HO5BDPLlBopcsabA5Ib/GQfOU6y8
CeDJK44JpGwE39vYhSEHCqJdRX8hdkLs949HbBrEZbuL6iybJ7EXiIMB/u6NawUEulud+oV8LU7g
Y43SuxJMb0HOLHMfdDCxFjTn+qPWX9DEXZ93gEyBOyfC/B5EE78Seaqh3K38Hc23TwP74pGIf6AA
eCFkDUfaXNYGmZU9hWO0jfGBcZ5g5rgu+hcAS1/zh97e7P4UgirzhfH3/6cNo78OEu0oEB62nPCy
ZW0CxxfkUtZJ5ntlf1/Bkqd53dJHzcVJAmU4OVyKMAREVBw0+mzA6C9DdB02mn4t9rr/jI6s7XZq
UUHyKWecbQ8RfLAz3lSS7ImUYXf0tF05iZezapk1SXd7Wwm22SXTYVQUIHb/oeOU5P4MaAgqElyw
Ge3kKVv/onsPxPx1iQyKmmkAZTgC4dk5lXyf0g0xaDlUZqTOWlW1tz6dVq47AT1fVgRQ0jQgrp22
3genUZXtPIIhdRoqUErCtFVsG8VR9pQ2RHC1krOBaRYfOPfGABhTUOvnDxt9TkBwtJVM202ZJBn9
KD+f6SFNAYIb1q/Oue436RAvGmePyLawG13Qsg+rQdBiCoKXNAc0MsZKgTjkaiMeRUlPcAXcVTNJ
ZKMetLmUenej5/r83noi62oOfkyXY7yZssyI3jriS3aJ6Syt0pL+rI8ij6EyRJ27b1Hb1sVoFbXo
/G1iQkvl161IS1SbPtXJT5D1pb8OlbqybquUDaXHQmce3TbWaptUCyqHkyq/yK05TQ+CpEKpp7F9
EopU1kORpsIhPbDPJ0xJTD217zaI8AP81X03ccO3hUPjNTWe/iPnWVlp9tkRPv/8aLCxZzvnm44h
lBhohEv6w1u3iRobLnytRsWbahgBbPlooI9IhybMn3proFstqHhbV722qRWW+48FJdzjQHSS/osu
2quLD6FEqzI0CfwCVxXMMh8I56Rzq9kWOtmXXTLNdPKegdwwHn/exXMwgq1RsL4Q4pjgMmEsVJbY
BOoytvnR6takpIwYFU+MgHJb0ZfR2alWy73MOsF0cqOi2AlwadP8tyfT+kFIe0P7yvfFqaaOGfsp
kQy6dGTMx3O9GZLEWgS3hqapyWdBoUD+UqjD9JVXtq253MzbSq+5A0jENuaN4I71m4nNz3w2H2eT
0EhTbbPQOwBFYj8kzThtKndNTe/UmxuyRePY5+jW8rc/khgGbUyz29okgK0Mu2CESJ3Ho/3/vhj+
n5vjTwdFfATZ5GgRgHxPUbB0ehrHQBN1QZb/gbRibB7qLTS033RgJNqbH9g36wL/R2X+VxNByUb1
bh+I1+FNjpqNOvRkhwon/tnQPZ8fujy0LrDrtAMw6mgwJZ66r51CmZoJhP/lyykgWpX84f51xkCn
AAdE3iBJ7wboQ/KELp8RR9nJge7Vnpky1UYT0nngQJtw7k+u0ziGrbZdNEbtZ/SBcXYM/Ri69LKX
89ta4FdT5gZyirsVwgi755Wo5m+R3xEmZ0qqaHMqi+etJeQggykBr2ArZB2nFHRcDZdveta4i2/1
MPzPlWWykVrkk5Zny9X61eEF1kxylEZNatq4Y43mBllQDVkvWz5QD52KMlbrNSXuj6Zt0CWP6tu0
kbEorfu42XKaaNaWtzK4bR0582ubEnNIR2GZhNyvJgVjReX9tXN0S3Bdsry+cjNZGL7xyxHHmO9J
bsgddRjXtqNCpGND0X2hhUPAorAdsZzl1ZnkRqdACNu0wkmY0Dkc+ZDpyINZz8qCTdQnBZMnriFf
ayfsri+DBy9xWwx+TD9SmwCa7Ach54sPSj/YmzyK0b3buFzM1F+l1l04Fi88ioKBesZfhbIgQCrX
keE5PCOF7lL4AZEvIB6ZRiFA2pg/YOxM9cRtWXXTyHFapr5zpQiCXV8jTkRlHqC3ZVvgjvhDfVIW
ePqHoXWBL8AL9Hr5JwrwneowCqMM+x0sSoDkwX5uHxhC8shGTaCwIA6eDnlo3r8LZAc4o8FxI6cm
P2I7ynYKfw3s8+H8WnkfTq6wgLJ8MM/mgAyKv3XK8RNJsiFpwcAJr6ZrR229v5+vlflEFscbDFG1
YLAD/AnzGL50dkX8jn5HamWXn42yJxEjgBF8EqagB7UJY4TLXaGI4ymo+DcNrDQXnfLnrxHTI6yF
HkKuw/qWCKfAijAffMUi+wlTsUI94qjI9o2MVfbfokq2OiSzeiEWOyjsgMRTdf40Oghc2tHgbLFi
XvVMoD3MrNgif9N1iPzlX6PnBAHDYvjqOZVrDwMrO0Qk3AFpwHif35Nrd6xT8EyO0C6kLyY0cR9k
eSvUkgwZE52SjYToZCH8oh+qoKQJq8KiHNms7LBuE/vrnJrQ6KjlOQ/5kNJr0p84ULZ4uZQkYO8L
XoNa0VrCLmIYSKYpkPFryLe2ZI/rpC6/y384+0ebd1n8TrTJ3u0dxsWg1vyiz/OO/0MyIcyL0jNc
m/rlgM7JEzhmO5VXfYg3rWuZyJw2SVSd898KF7fv4q2cwN395s5JaE3q0wKY+xxXjlkNyJKb24W7
pEcygvx3JkmvJYXRUWuQEkM0T5bXpEOZNgtnJ9zqZVajvHwMY3j6+OjzaT7ysMTOSGDSLWk+xNhD
Ncapcg96zqcGQIWIT7RyZbK2Pvdb8AUUBVtxHY8B9I8fW+ZF6yxQ/v9RKGKNB+uXo7MfIVw3+q6u
CkIvxkIClkGfVDkPB/4mVPQztfuWLUQB8fhdGhsbZvNMAySAjXeyqgzZ7b+9PG6BMtLRZSn2wuF7
pL0TC0Wmko0umuidECD7gUmCEpxbDLj2TdVe3XrjD2mZqdmrulGEvqcBB/3S/v8WfffnD3dkej/H
Mm5r+6xBY8lPh3w5yOgg9Bk1DmI6Hf+NVDtZZFmdDg+F/gUjaeoK3S/O2HrcEB3RKPWjNwXe3dX3
qhxK3XsssHU6+lmcZTP/1rtcnKpHtSk72s8oGufZ9ih5KOIYqJEr+/eLp6gJq+ISc+l/v2ZsF0S7
/XOLGHoRMHI8DDxDYgzSBpDPZlFatODbKccVbfoywq4Xsuy5MdKCFQeDOg6w/fRKvmIOTEVBvVuU
+pAuwOQdNBvrSmXwaQFEwcKJvPKLsE1EUeZtocSFGjSgRj9COTr7C111aKwBUvg+5K909orCwuVD
LKfqGHaa6fK79Se1oYLBoJSBgDPnw3ri5uc5DMUxv41rgcNQN9v+Jrv1N4tqyIhdv86z/5vPwPYi
HXRmwOzG5SUqoulVlv/KaVDIOJXxyYcSu6G2n1CnSwoEy2/Id23ErLOfR8xwHFvQvqwVUGz8NTOR
wArro2kfJcKHTtnKF0BEMkqZaKFexZoaOhNhFURRnjU2kAvvh5I6ZyHkPbU8rMynxXrLu5n2ijAg
KgbHl/HhQVlSgYf/q7rY4m2Vd9zeMo6FbbNypinNCk3aJUGVaNDVR69nQSrn54CpBmjgvtNh4nl9
KavBMTj4ThtLwu4uywcu00PTRzzA/VfEQIOWgEa3gF+EyjSiin7k95kC4Agd4E/e4WzcLbGV6zkh
a7j7vD1pPF/CT308cvqqcAcqkIMX0Oz5dnDxg52B4qcjRqYUmzv+6LcICOjNqajUrjYGG5++bibI
jwOdAvUcUE3A2owrHr2mE1NfEqgflKhfzrIF4UEesi5KvmTHtLozwb3k9/6Enr8HiNTAC4RiNUzF
4OPqjpnZLoF/xaFcy23mKJfPmnA5KB9CotOi/wIyt/8aOTHu8X1SmoXdi8aDjXAuBKcDynDhXGkq
tCv3IseJkYvvw22xcQEfBlvJYwWAp0Crxg7uzRpFvBa46uVWAHEhA76MLcRTQdzoVENoRSsxtFNd
WPAzMcWFZaU6ZRf4NtjyuWjpr+Spl9VwKYdJgYOnD/ZlhfF10CAdc/VRzC0eD3QBi7IqnH4QaWGp
vczO+PE9FYluUvzsWsJV3dW41YAulj0E+Nu9spEIuXjErQG355raXhZ29/56L6hZvwGprv2g+HeW
PcV/zGdXNEZmd/zSAsGNiiwfWzOl6wqL3DmCtCW1cSOYh49hoD60pmIi8s8h8BPEqvJatVcDRnkY
0bTx/TRTrsKERtxS8Hm3RY7NXiAoLj72TjR0FBm7GXABIQC1VHbmRWOFe377BnbVy5MfQybgVP2n
BatBR5Rv/SN4LcfIaU+c7CrTjV8uke9Nif/T2zcC0sDbASel14g10EPud2+I1JfthvbM2MTLvgYK
/WRZMLUMBDJlfylnuXZKjhxybYOp2Gpa+T5BoS0EUnbmIX88+GKwdgC2YBDb2XWn5Ut9gE5dUa7o
JhgSZqoIMkOLAc+18R7zXbyfTYW2H5KuuttRYCP4g8NhXeRgxOTJPOTNJuQIUZSgFRgK61VMqoc/
TV1DUErAz8UgW4nwmZ4+gekQ55tNh87f5rkg6d2Qh+S5EJsWpRS9LH0uAdzMkwy+idQXAB+SA746
Y4naKoBUbS5JlfHIUlt2mwHWlEkgPbGGjU0yU6UuBrqAI+O3vE7dZNExjGdkYTRiyS7iM+K27i5R
/gHYxQ7kSpQEe7IJOnzxDvOo7mhuqvJMdE9tLnKgshGIMbaSMVyOU9omD55Lr3eh9Cp/esL06+lI
aC7mPEWjFiXDWkp7VSqYMNGmNfKO8s3t++3DKYvE8LoPdzUz7g4qz77LOMyUOTg3z/6aCo8xkfqn
4WNumTn5W8VOZHFSogd6tuNdai4++HqCQ27yGCM/wIMdgtKQ/22BPcClctpepzMHnmiOv48HUJGY
6zAPVonvN3X34HX3WOrb+NSx5Zx8alhiY40fPX6AgBf/eb2AhF5bazM+8PrV97UcbDuxhiMnq6iV
KraWRcb2GwgXZy/N2wyd5PrUlAbvdmfUHbugCzSaKKIYGlnZoxM0iC4fha6lLHv46AGGpsRY/Aes
WUhispDjLvm/wx3Xhj1GD7hIQ66zuKqlIiXKgomNzQxaVkqvA5+YjK1Lovgy2+8hKP+xqsH20chA
mHLFk9Mc5BrZWbPO/MAIBlmbK9T7T6lDcB4Hs3+9+05D0OfZ4rONu4MgWHKJv872mccaIWsT5lY3
xqqK0bcn3+zcA0L1MNHzBnNtaDSa4b+E+0Suu/x5tHjovFn7TSskcoyP2IgIvr6y9AJAVIzP/7Ar
WiBfeFTHCivT3Ck/ztvxpxOR2lCwElF4d8YRA4/jyi8UqucG9SS1zPBT+Tc4Ia6QPcVva7itB6Yh
5Tvbde/XWaUFZbqmjIGjiipkOzn/0XmzNljQQCC4uYgG9sKbn+fYcSdvML9xBaPVr2+BevNw19Dm
e1+P4AhD/wdu049OLWusrBU5yOYiRQkFTpm/2yhjnaGjQY8l5dR6/vmNoms49Dd4z1TL/MWjcF0S
2bavJ8hlQZ9PNXegL5dI6GU5OFcf0Rwyr7vOdA3xGTJsrX/Hz7qTCHQsXkyGJ5JzcwqT56rT55xO
dKVU0soelpGwJpdvVIYB89m9J9jjYFyblhh39NH4LnkblosnB2S2V0wyx134iGTxc3R67c4Xg3kz
JB1ilRdzi37NTybvcixAasPqlJOF+7IO6+hG7xzcU1pVJbsZbTt8zhfeJmT3T5JxhXZVNlm0vZXh
AR4AihRSSOqgEpVbHMcaDBHb33VacdsJ+TXF3NV19YAPz97dVB/pNWzJQUhp1mQYRorcmpx6BtFn
lhN8D1ITfqA61O3LLA9BEgac6A92viZHXGM76r+KDy7OvLRR7BgNaztndm90Tcfi3VHwV1x6lUyV
9fKkyFo36xaq3TKikCqh+L9ejFuar7KtCeEM/s9dnmGLrl22CWClyDqHaSpCtqjRhFkbJikfCN3Z
Gr5hjNKQvY1/GXeYmCJAdHncf+/71UNcAnESy6PoknjS30RG0Eq2kaC4NjEeDLOAQB+f/0LRK5/+
cOffRYaiB45Y1aD3bAQPsEDw9FWh4mdwwx9IsGzCpKYtKiUiTbEE7gWfpWovnfC2rVtx1QAzhE5r
ke8Rsz8qQnd8IWgi3tWw/Pz4LXw4jluQfO+Ri0cxNHyFN2QmTcH0DlyHGTStizBbApbDvtmqTtaG
gzYWQVkYu9qxZisIrfKXQE9IrOj/3eEG6TPu9vYrP+fOPAwcLa4OQD6pYWUsiACfjyHP2ETkoz66
VilBrzNhOiB9y19QJ4O4jIKTst16V6fEoSX7H9/+xy7uUBNqLpyL/nnAxChNqiqKhbF5x+u/TCqz
CISBl9zJ7IgFSjkOt1GtcQPCcUkR/HnnQX2f/PoRm/56nIvd3uddBy2Zrjt+xYBYVcEKUBzfWpJ6
t2n1spD0LLyNg/nhK5RJaVpieDhwS9VX7DHNB2+kqPQW26vGB/cwJF1rDfdB7HRs+QRSlClN7X2f
ganMSl6cifwzdvhK0xIjHVXrqmGIndBIa9FVA/C2sIViKTuJZJ0aioiy0WqDo+Da4MClIr8WVN7W
z1xcXFYRs33nbJZWq9vn37ccnvXV5Q9OESjdgewqzjed7CNoyJst7O/6TfP01Jxx5PM4/RxKCkJ0
3eAAsur8V5CY9crLO8n+myAAexVQLq2xgg/+RF6GJGuVSwU2YHacz/UlUQTYjQd9W4ArWezqY3gA
Hx0wYC6XRoOE0/XELniPA9ErJpZcNCm1+HQe0olpXanAmQ66hRvhBC146uwW3AhE1ksxTzLoSIyS
GcP5iBnQv4otNVK3uL9AIY3Vbb36qy0FJCKQ/TlUpDpLNtCrc9keneJAhQmXWpnIEUpHLxfjEwff
FD47zi874RIow4qbiEI7SiEULjIH81trIC7QZLNScTR8Joi5j0t+wg4KUXYZ6yYBfVDSk6WwqM/U
Zh/nKlDNY6tlMIxUB1aXyBlgAHaQBWDb4GGwLYkGYoIr+IDgdI0QqVolHgUK843kgWqOMUyWIZIO
BZTKqambbC6HIJUKd02X62e6CU3EMuz2k/ZBz0MWjsZ0i4MvrEOHUCYbnIUyr7spUWY58haSQNqA
TSiOOtET4LZi5Cx59tZ5ijB6G7Ny+06pw0O4gNESBzQtUFQrBmhuhB/LV7lDffIjkWHoJZKRG/0M
MJ/pr3PIV9r1Lqt7KSKIj86AqLvmYJqFnmQPDnx2ZSnODamVvjqyywMa7TwNiOEl3bcLGLsc9CKJ
RbXprSNCtuUcVn0reRXYX9cbUxZgmcLnqGmZwGcDltip4tiirfrPO8CqQLQmm5NxIeiFwz0/0xWu
NI8Ef2Z/7f9UTBsFZCAKzl61GRNEonvt/O4q2kAU/5K1ZJYOSVJXb0++WOrGsv8Lb2twkniW3n+F
ykXQw6zIjdhtUV5npUTEsvjlN/WsVlQxbHs5jEPasKDfEEmu3Tpu0cuXHTa0n79Eu6U/XYBRKhZq
eskl/DtzcfuGZevXG6pUZGBWoudocpbOpD0bdTaLPzzqH7JVj3GTJDud+pw0LR0aUA8nrW5MN/vP
0OnNsbc+f7P9vR2EIPV/k42rEONtkQrkrrwcZ1kxmD+d3abRzrwEU6M5Xhs0swLUWP3aVcdoyyz9
oeXZsbVtYMKjFOr/GxUvQBZ4u+tWYRu/Y2l5MxhNGu9vAMjwhvGtKFbdsXHPQ+DshWzWo/dcigRE
rPJXVIGKq6hvBLTUyOEViOQFNBNxfT4VdVFPR65CcGgHkK1gAXU8UgwSgXLIbh2SDqtPJITdxmIL
mCfPvbUHH/rigvCT6QlYe2af8uKVqa8c2S0eGqRrWkZX1D8PU6yz51aPjFEGtT2YhUGKAlRO7Rrj
n62dd8ATTSZYFwsi6O1mm7bIxNF3tgha0SyzkHgeZIPK/hGTmMEUp3covEiNS9WFVviwUU7Km5Ws
baq+pHPnWHWIo8aPIizCN7o08Fr0V0CUnD3NsEWFG6N+smlRvjALmSq2IyqAO1/RZ0j2s2EiYgt2
7Q+cgPdhkbkgy0nTNuGhLiMje3pVdsUuPca7Swahhog8RMArMRmTcCB2XSoSQIupcCsJwZsgZZau
CvLxxyFOov6Ji/aY8hzXv7QDGRGQJItYXiT2xik9T2dlaQUVWuLKj9DCdrjdZIqJ6T0AlQzAPdDc
L3D2R81wjTQrDgAhYs+dtbI939x8amzb+3yYYdA82vRX1wx8cY6r+5QQ1Ven4MyDj9JMOmD29z6W
9dHH9S/AbZjjxF5LH1YhtegcMr2f3QhzmC0eDvml+y0sB2NRmVWQUlAx9JSMW1w8O0r/LR2ZAsm5
EZoQZ08paQHxjUQ21aSCKzsGQMnBNPoUQ5ocmTZGktWZegwzJtt+KKb6NHDRamwjApFhW+xxCmfL
jpNdbPe427Oi7DOTzo+Hgew+saRCkaoGFu2FACZ/UPr3Xuft2DVOGmYbIEWePgqVGOCCH/VoH+5I
150EfA1pLtXSdKLzq1QNGiC+vA1fG9xqphief/NbUQlCIBAkqzvojJHmz1jTxMnCWmNmvjDiTJIO
pb0dbF4Vij8DYsVvi00w8yp66cmOcSj1lRJISuwuneATppA9MUgPUpmK6cdwwc0Y+ausKnUIsvi/
c6TBo1ad+/527m4GzG7sK8HA5QIzjGmmY522r6mrca9HcT2QKB7SSBSqkn+nD1WRQYngOiRJlAk7
9QY+ku0SBdJ3fzrUvFuCZ0yFMLd7rUW7tUzhuw5ZdHTorIy0NlFKrQ9mS+zZbQO+4/dxEi0GCIZN
V6KF3t48Q4JR0UDNWYRQb3HQyS5ZFI70GZGRqxwXOnAJp5gfZCrd3Di84er/MtULLXeyFXvzq18m
/SEzYT5Al6K4GiNztrfW1j4LTMsUkzeC+kva8VBuzZ5dETdU1wqG2eDDl/Cy6/6JrLPWg8X67t7Q
i/ldekyQhqDxpOu5a6ugj9I33X4ieVi7+Hp39e0VOCjk6P8ttcjeh8GfjN/8ldwZFhehfDi2ig4z
Kkxbz2E67tGH5VD6EwAm0HNWic2K1a5gxe7ZmmjQ41OLCN8VZSDzeR54hHQ7hBLZSVkTf5ZbyIsl
O8yRiUZbdjAxoI8atWcAs/mkwD3+ZC+ch/5krvRqEjB6mL29Go5PA46xUdRxwGNhKOADh8OmI9LD
KK0Q+aAQSsyXjk5z0A53xuaaD2ZfWpNZMvUgEJAhHI/bEz+A1Lyy0OLrkVzRBAVui/lthJYV1ckv
oVvHFJr/a6bgon7tcfmRBCfQXIzrMllX9OX7yzEhkoTiQ9hKwzb78OciJ1xSHgyr63hZ8MSt4h10
I7JCiHh4fx0TkEexdqoy6SlZrBHD0E7CJbPQQcgOeIR8943NGXgb+BzgQJZLiDZE8ASrr/1nnxby
l2E6P/tHlEsi7aCzrodFFSDb3Gyfbl3CEYBcjEYyJGZ2tWNwXaz/WkSm14pdR5Ym0nL4Xwu0Ccq2
cHf+6DlMfRNfpOm9v3vleRG71NGW+JAC/w30p5UYCuVi1pmOrqUL7rudDFJDB2KIF4n9ktIorGWv
JvPDK1wtVN9H9piJZXdOV+R9eF8em1dsxvF9I7RXyOzDiBAgf2WA6kRuZSJWuKcdydSXD2CTR8lW
3GJlKzdE71faWVVVTR8xfkUu94QPDEBr9607U7H/drN8+bvrcbgtXD5iruUV6DBNeN9Eq0f3D7NF
HOwJFb+s3exu3kBumfIneNxbl6Se4keZkWH2/ByijV3YpWab447awUIq4dLUM7Y3o5qpp66/8nWJ
UlIGJNzcgt34Ax6lFlLbho+jjh7Q2WC1gYV0YG1vepEDdfmDPv0F1VAe30aiW0xFz0GdZEaU0qZv
MaIS/Fb22Z1SWHYTIg/NHmiaZicSpdgq4F0UguenozU5Qs84xXrVR/cma8RUOXwQWY9v2yRl4SL7
PA/bzwkGmUMhH+LzrqY3Nh8Pug+KhTl7OKd4hYAEiA/JFCdCGntpviTtz5sHCVxC1rEoTaT4GV31
NyeFL7iQw0YiiOz8+4mbkr+2Iq9zgO9RV64mS8etKiTKr07/WP0XeAh7VORzChyM/h3FZaDBp9u3
LmTCtiOL8vjwlMZ676u7JmA+E2Kajc50EhJpF8YYg7tPiFot566hMeJVsi116Q9LZxUELxxdiCNj
CuMlGP+Mekr7U/q5YL0+NySx/rHBXukGJjUA7XVTBordD149dM6T03OH46reG5qmt8yZrb78ai7v
5oYFWpDjD3vXw04EVj1kC5EcrGXMYOJURkg6o6Q8nUlNeW5l8TDiBlZr9vz5oTBjg4LLAzr1oNXA
hqhrA/O3fEIaS6mR9Ake63IQ0Wubb7U22NpX51A9UvAcQKGdQvWcrfn3ib26Bwipt5/3F4REgj5Y
Hqa0EHglYR7naEDPvT85GWCmfCIaBk2NpxzI4LX1govJr4CjFuc3sdeh9PQWTIHJ5eClQ53JJxOE
VEfbAEOgYLqYa2gaaqNwvR0FMM1Bmf2nIWFiQ9lI0NV2O/wLY2k4RHzTgdgecS4N0rggX4oSCyLJ
7r0jbdv8VgmN5xG0YwnhtCxV65PavfXj22vAfppf6r+h1wa2ewA/9+gD98IS2zX1sMTdhqMHoFIb
DtwRNISZIzbllTPASMDhiWovWeJjrZfty3RkYNM31SiM8OcITsesY9YUWJCGpNvJFVvIuTCd7/Te
bALk/aaCNhJXh4RQQhBp8rhyjwvzJs0B0CkTym8a1bmeN5vrrbyC3U6+Hn/v+p9uN4Pipq9P0kop
TRfFYDVZhkpG7b0Jlu7D6CUqHCpkG2SXJn48FWdZXr+pJbn5QGXYkzLTvxcenIeSlCf/M2aiKGwR
joLHAqmFhDnSA1Mdprc+AlruXg6EPzee+aTG2JfMJo8e+OS5qxY5C5aJsAFP17RJSIF0sKCkXVkW
IirH/YM/BpchNGstyVLX7mBBbcOAOXI1fRYll6CqA0pDP0ZtdednSINoWYHt1y++H38lSE2LmKg3
FMgCedx/BPpyahcEs8vOUa+2pjAuLC4AGWnP+J4XZ5k//T/XX1G+n2W7cZUglKJJWfdIF1vYXjGl
39AfU4eiHj9AQ3lI+Qot0IfCl8QoKCjNvHeSuQ2NMyy2/56wD9XxLWBNVMaffJXQyOXg/M27dimg
Kg2Hc72jTpaAduxvO4DwJjzjU105zCjsvpFzDzW9rKL/TSq3fsLoO5L0MLB653nGDoozc2+fh1PU
VUHpFh4Fft5ANlicQACOWYrJbT7FqJHB5ORkT/1NZCAQh3yD/DVYIUz7TiTAwJDQ0dIz/hf1HWnF
VtU/K6SfF6TLeeVb278n+pBAz+OzMm178ytABoPXE/g1EkSOlh+afJiAA8jnaugu/JsRH9/p7/wV
ZsbZBqCBqpDMEhWJSzBAVgxShvKWTxtA1I95Q2y/F33gnv7G9G/TRCyQLJHi00dhaykgYPkTiwJO
tN4zwplRjt22FwsLB11qB8SK2tKKtRNLPEphbYqKulN8iavvkbD0DKQCrPB7THsjk0+k6KF/gVtv
DlcZK/NoC/OUbYCRb6Hyn2/vRS70IIcmIox9jxx0Ed7N8dVHlqhMO49FU5qGegx/TlbIwCT6VDEG
zf4QHISJcMTINOoXk3N/BPcLFU4vmatbRWg8DemPLUmBuq59MCAqYbyBrAjVD2CddT1RbFMCIioN
BwGp7LIxins+PdV8KqoNKT7v9ptqMWo0oPW+1beppJjmIjc2pOIGLwnfjrYuzQjOBFYrd42su8pH
KjsPfIg36KxxjCPQaJtHroLhz+3i5ZqnPQMKTvcqX4HxIx5vIWUPE25BKgE/9xQu2lNkjN26haiZ
7CJDEePM4iVxPggQzP7BZjr/5qFJpWZnBo9yOjT1+gA19VKWysoPEirNHWGn+qznKMwBPJaLjb1J
pVDyxd5yl1prcy/boRrVJy9bUVH0qS71qO2dFIjdzvR4A+ycNsewJfSe9vQJORgHcRJD1fG7iB+H
b0/LExzFGkatP08QJqEoutDugrEUmt0RWfT4ZMUyet972r0FukU0aCkHIiS7jbIiv/XRYFT5gDy+
KVnuDVTIzsSb54MY7GyDAnvXiEeWuhjBYroqlaPQPwDEon88VMVbQ6G1TihSUliqs+KQIhqcdSLH
ArxY/fAmyv26ZJVXRAHFB1QNsFP1ZoYbj8YBQZR1aD8j38mtxZ4Apr2TwcDPv3jOSFbYycksaeoI
RS2269BatkYz9ShnZa0j5UEqc5m4nf8cE9YB8bfUEPqAzHd/selZGElYJvJNjT3qAjLBWZMtqcmw
/fMrsM7W1dkuUUZiuTCcSEHbGKN0k4ZKGpmMZZDdjUjK10t3DmYVe26H9qdy/V+Prg8Z2VhZGf7c
DhYp38gisQyCLCLynrphQWMI1ovadCuh0dO1GJgPa5QoiISMr9LFgCzBY2tsNbHujEouhxZBy2f7
/Umnm0RpDPFcK01StECi/m3NuqdV6ff48I1Xwa/rmjQ4XupFycR0Vj/3c6hKQEN99JF8/it3wbel
/9yaIcro0pTHk3oqGCqJc5FmdgQ0NQNxnalfGAnzmA+wl+ZaAPT0wUWV6Fc3PL4c29lLcZvuOmzL
+ITFde8CKcjChGecJTcVsfvxNgDlhp0CABWy6iVoNvmrMEb7Bcr2pON9fhgazEviIdq83q/Q1RzN
7V4D976zSm1ccmSY6FloVPbl9WD7Pn+sJf+83cEbUHjBqBVyP2AWJ8q1uSHtQfXc7nmKsYWYxt6m
Md4ZEEM6u+rn+shz7kpd2Wq+Nm0CCqguxl/YTQiXtFnFlUDXMTC0LJgEr69wSdgFghdpn7Nz+jqJ
gPTlFxt2gtODP/TS5eF7apncHbeXE01feKx1rANfjIyFysBkfpnZ8K7ikzUHGaU8coYLTQmZQebD
Qsvd+GYu11aRexUN11ZSFBFnAVqPSBk5a9htN0lA/CsEW0ZrSjJukFuGzj0GfY5QjKAisYMYG1Dv
EDdpKmjJvmnyzwzG52C3r4LGbsrtSFkGzRrDYHAp0HFW6xV+MZrV635OAe34QWjA3hCNAiOHT3s1
fkjomZgdx36s730LaE2pjvUjk14MAIs6owqNwOMFkigRDLsX73p/5AqKDF5nquTXgndA7E4qdP4a
NtI2VfSGvFChaBaOv/xsDaGzYStes8haIWdl8wVZGK0wAQNexQelkXlPE+2N6kg816VCDX96LTcQ
u4J84XeeCOD6JXWYkUHoj5ym20kKfxIlxcFkLBYvH67rC8IVCe0nZeWaImMVgZ+0X5aA1EqXOGIR
r6guHKpsV6VAlis/gVrpS0sMj3+J8x+wLWdV+pIthW/zpASoldZbv4BszrXzS8WhL8+1vQo7vj9K
aKIyyZ/GkjrG8GBizdxx3YXmgrbjbBe2Kch2yS1Qc5NDF/IVQtqfkoI39t+PQR2QmDUz4sD2Z6xr
snRlJG3SHnrozCadStYEVGQ2tN4YjV+X4WxuvNQuAX873kQTnIjmuXSjlZVIuYge33EcjphSqpMZ
Xfm7MIeHW4x04NnTNdaCXQaTpK3ClQAvarQP2DpT3u5c9nYjPtjgisEwyc2bGEffSuk0qt79I7a7
qyWvoRG5VeokEN4xBYhbczn0Etiu8LQnNrZjr0IAN8dlzAyhxwK78uY8EWWwhZ9BXskvvh0Enuc6
wrViiMNMgo+9rTwtzKG+jIuphkl0xNEYOvrYQebfcjASrt3wzG7gfZcD4fw/TBIDTa2fouycoNPb
15TGUEqp33DVMThgOEHlYBUZ+jxp0MqYiP2+xRJcdVOKmwMGNzJgzBXzcBFHUR8hWJg6nVNx22Wg
5axA6xr29TFfpBqjOVQ8W/3N07/T3V6MFDAvfXa2XYTwi5X7/BBBD1TNhSs9Im2IaZKjo/TLky6D
qQ2y7iZziaCJIXQXEbbN3Rfw6cOl/fpUzOR//gEW6RoK4AEAGDiCsKoe8waCVwibcBxeAJXJ8rI2
eua4HiP2BFRGFEji5YwoXbvSLpotlAOV2DSvs6JAHyE9vh/kDfMci4dcq35++6qkfc5EuZaiiVI3
bmrOictshd+77mBK4Pvo64Jf0iS2JV58W44rrXR15l9gCTM1Bf9k0KhM6H5N6rEI8c8qE4fzk423
hAe7CQTxn50KcokC8kueNeR88YXXds0rwRfIhjlafS4j6wNWErIoYMRp25BnX/iUlfEioyDZzozm
VsVC76VjzF/UGBZNsOo+CToKS4pSJpha4qkTzfgFjWnkeARndT9qv6xoulPzT9GyL8IMDrtygMlM
CU5z8lVWxEEp+464f0jg9xs/I2UJGZsgq1K5wmR5bxEYMmNDRdQJZK+qVqrkyIpbzKsTYGSXvQKN
aaFoDdhQ5d3y3keL08eegUIU6blgzz5iHIxh0lAixgZWlxapjS2KhoZMAmTwgpXCAXodQPOwD+ci
uwSJ5dHXqsaX2x7sHHH5J8hgTFiVWauqefd1KB9qYKabhOHZDfVRpgYQV63ivhXkBCxIxZDFIWDG
OBK5UH9PLn0EBDu7Ahbhf4zqXFe7BH9XSBOYuvcgCLEKEhHAwaFhcBmM4DVnIVenvLv0NOEQ7IxA
oHAqodjbinmOjfB4WN7kW6+3h5J9LXst8UNVdUS9DwmmCYXxHwbSjOLXNdoXu3hInziwoUPUyc8Y
9bl3w1uyCljt2BzSjpdHlHZE94HRIGbD5c5d7QbicJukwgZx5tUKtJu+GaXxZ92erJ+TJ/WdtkOo
FEtb8PLCfQgKsz4IpCwY3WjWg8w12dBmyD0BJEwrnOqOM3Gjp7qwDwlbnGkA3mblCi4tFO76TaqW
6WB5JQNJzC3gAaoNZmfET3RoonFl2EPXKpEt5xKzu0ORTOPunWIxCMIJF3r7eQZAjt+SfhP7Q+6g
lU6UWRxG+9gUM2UxrY3sPWV6mzZO5B6MUWqtPZ9B+GulycpZIku/rbKVUf7ZWaJRsHOZvUV480B2
SVeZMiHS+jKPV6JqIYrdmuuuJw9cIC2qM6Qc5ShXMFs6AOYLS0vIcVRB+pEqTDM/UkwaPGDYsbO5
d/ia9K+PQgRd9tLbs4MVR0mtNaNko5HDN0yEUnHnvnvvVfvJc0KLM3wWSZ8sfavzquzkxXYfgkwF
oK313M1m3jQYRvNcivoLpRtLs3o8feCbs3kE+USW3wS/i9dqFwuryRHpwrejDmy96Hxfcob0aN5R
YOAJc71JXSDIaAG5y9fWDG20EA4T4WKTsFDNI9lpenZ9YoCzeA0G5MUvohmIc/EyyWOAIjuin8q2
cwBnsNUD2elzPiHTKTRKsO9LDiXhk94vqpz+mkvOsfhyhEaEtA6h1aA+/MSEzJtQ6i79Sw5O1/0U
ggAFSOBV272tESoxjm+zuU9WrkYlkX9PbUnsB2mBkv55AGMjwmqWNempQwhEQi69icY+nz9zA3eA
xki2SPoa5qS1pm0j1jNxOBXxlH786ImHnLLjy3X0o/UsKfN9RtkbHnPmb8AfLwGuQNapPyXKFoFP
/yqZmLtEcrilJcjalZCb7oeDY/QTKA9rLRs1qu2f16CWAeDuxb/AYVcd1mbIpi/cK4XQc12CVSy9
KpbnsjJhLmdvbu4jYD8Xe/hJ5S2lDrBaNWRPB0GQX1wZfpmyEbcDAOdib3tPHkgitH+ROAE/AmIs
MVZ2NJFRy8EmysUU42wi4HbpbHwAEw8pWvlRwTbsMRGjeyKiAjRKJGMfmqhBBe0leexAWuYEFU65
q3GJORFJ5E4GMe5WnJy8d944kJGOtUDoT4aqd75YQWgTBtW85cl6XHbR7hb4Hcj0OChokSvOUZqy
DE/v9zEa6OgyFrQoZR2XiQcfNZjiVMpz6pD0nFxSCCp0OmB4/Ap6iF13cT0eKPRSGP5F7ysR+zFw
+ey2/Jv/Kv5ZCT/Di87Sd+bAbFBl6PBca9giKn0sDi9ShLVfa0HWtjwUmblSYeu6nO2Mt4xqY8uk
r8cfa3WtcKGuMAzgS2MbZrlepaBRK4VqLVTg7g+bT25JZ7BXaEiEQYsh8njaOSuAIMdrnsMBMPuj
2vcDitVwfB4cN1Fg28rI9ZdRA3jSqPP5e5qs/Nl+jMmNYU37B/u1N0vK145GvWzJN0kkQExWIni8
BeI7+osQY3ZCajQdFyufVVhFPu25JhWyrQqUVCcydrqhB1WXbGs9NpCMflytXuadwgxW0MHWPtLl
Oz3DWpoyHg1uwBAUutXlpzZKh1HfWV33gQ2V3pU0ssvy/GiohFZ/3lIFIqde7kPoi69PN7sqAjij
CYLYQn7hxkHriGsH385U8okmXMnTIi71kHD7hONvoSw6a7ho650l4vwv+9AiIJlgy+YSwSLSgtqX
XDexW6/JWJT/nu1ulHHQJeXO3cBpM7auqBlTIBZXokP65Zs8/BFxo5f3cZJ4sAexk3dmMtlFnhOQ
BljW677J9X3kh7KvyJgH8tWrehXWtfjObnxQwblNibolzwX+pBSBliETHI5dqONmO/CvwHIhfIyv
egoL5maodlyUYB+ngQwHU0IfGNUH/bcnYM34DmLEIbSSd9o6QCvMYm9/QE4gPXauXniA1PGYtK0L
q66QxWBfrdBsuBYY0EM5CauBbHognTkgRaPPQ8u7eD5ul8209lTcFqyzsHvXxV8cfrhI3lhDbYU2
fEwGkA7m7y/KR6l9UmKSTiEWISL9trp3I1dnd3Ga56L/DwOXtFIO9zl6NtF+/+CY+WM4n0V7PDv1
U98j3VfFj14AHDWvWo/z5QgiijqG7aITQdjLNn+mBHTsM76ccSKU4iL3SYgEJKBtpLRnrpAiHjZe
ou1IbRliQYk6TH9GRH6gf3cDSQ2RYlsiU3LrZefzegnFtD2pvfpj7c9LGteAEXhFY9SmR8VM1JG9
GEO/9uZgVlMKETuMqSW6KMrWq1/iMqOvE9ab7CQ4rqeRCs/1+WP2Oju/9Mp+laeRd+macfIaYUfb
6ynBEFeKjl76+w+L0zz0RfvJd+n6m8Ysiq7kIKj+0FU7XUB6jQhMof0C618o/r6aiq8U7xC82Owh
iZIPa6QSRP5jkQha+U7c9nBCdqaYjkhWMECdYjIElPc+Y/s4IfFXacEcec76fqT/M5iwS4G7Y7Gm
LMcq23TvLgwFctpfU4+L9kYgHxnJmAs9HB775jxIml8C8ZdQj8obX7RLl1mOL3XZJdRWTTeaU4Pi
I1IH3RkbQ9clJgbb++OkSHO+X4jclT5LdSEhlcb9GAkeXG0sln9or7Egz6leP1/SPc3TG2CbtZOm
mIpmNWwKax0FIaCPzwPmX6vHQNiVBiasu1OW5SHfi0Zm87WKWGp/OcmiPDJIcIuZvZMg6Rx2TstI
ZU8C8J65rGAqHDljWKi4GLJS9sV3dBshaLpAFwT/u6Q4jaOwutU1pE1uPdsyzKJWQVB+76vfKPU/
62mpVM5Aaeff4bdPY2aaDUiFv1irzHKwgThDiBfoeJQIYSVbVbnflEN9FwuN70HhFc10kxVmXyVL
lf9LZDMXo3VoOJN7BLem7Ka/6CoJNH6mTMsU/YklXgAziUPOopFBVhqFURqFO3Pbp6Dz3oKSCYPu
5iy+GszRfcoWhtTPkPLHWsjVrO3RALRsybCBS8qMG6RrLrGB7P2bcevYOHWW+B6rafsCkRQKJuI8
ms5NjepKzncEk/biTPgDyvg43BaDWv9IoJhAqF0DdejfObQ8NzOMhaH2iqJgsGiZk5bxhoqcCVq/
QroqKdbisII+4Mzi/XTfeV+3oKaUc/h9S/ZL6pfN2D7th9GaVevs4D1+9qtjp3kAV8yfAXlWI7yQ
lkae++FMt2rC5HLu4XTDKVW0YzoAzwLQiLdVO0qDkcjChFuPsZXYcjdxtPSsGS6WVaS9AifDiOz5
EZQNNHb+uzDDrH/kCOjuMnnlWQ+JnNmnAQr9owTPe1Mfxej89RTBSKZFWvwC0myKmNxztDXBVuOj
4sikAUmSrlbLh5pSB4MatD2YOvl4lMDGqDO6AGAK0jcQdYMOMYbn2ucIs00yVBs56LkhYzD66hz4
3n8fVLRXMRJA7pqT7uy0JiWokwzQI633tXOERaE3DUCZtOFjXMsLzHv4xs0oG+OEwDj5ENg4fIoM
65apkW/XJNHTgyEMMX7kIXWSisyWSJRxte6ZOMNhKLhKRNDsVk3Yw4IPYvGMOPB53mxgZaNhvTk0
xgHBvNrkMFFpI6MCa10kF51Nvp6ET51oKfAMFQfkNyoBHKAoyr9JC5XA/1CRYod8y/6+5OIgQZA7
UXgbw7XSBlr5DY39LKBOeye8zuSw9nY8kmA+N5AgnUKmyvhqsZ8dJ0EUZbNDMagecxrlZc6iM5QQ
5f9k2OJsFFY1KCiHQJbJvgdU4u6DL+dPdAns5jsLsoxLYouQ9fhzJEPPFJlteyzwsNpZxHA376UV
1U+wYFHliBhDi1+A3v3hLgIuG880mMfbf9YZFn5tXLVnT5pDvjkpSgAFlxNCttWp19PDoxVFrGOg
f6S0FEM/JsjEjNHVaFLEJRkjJuK978YPHIETYFo3/a/6qil2pbWpsIfiHxOzd8Ecuj+OMrXADkUX
lf4yeGg0ZKAMZb1vD0oBzO3VRMVtQSPcVYht9hHme1afVWdbze+4lMowd5m9yg35OCCspUINc8yE
1L4wM3dcB3h9dN5vx49h1LWsszT2CHnxdoeWGUPaRd61T8hLelvK+zrtprnucTnL35c5YtWRo2kC
eSjRedq1opMxs6PACr0vKqM8HpyBBeP4NaH5gcE8L9coo6saex0C8BkLoA12dodyrHkUmxYsQrNB
/XYj/Vl7VVrBrHwHqnLZghWxvk3ICKhlKCnS1d7FPnC8BABQH4pM3vXl9DMQrcI/XKT47ELxFYlX
TcJzQ7KbWLmZeS2+BthY/hheAiGVAKhfyPAUTVBFlrU0g3Da4N37ZAmaCX+q5yx0TbLxZPj1gdBx
VUsazgHo8vFk7Ql5EuOF2EtazuQ5lr8pIv6HSTptvgBVCvMB4ybR0/iojEkSeisL5AQh9yc4kXar
PGVSaFZXkCJ9k/lHhDKRl/ti2CV8VsqIn0R82Rw6HBsLGdQ0MeHgv2hOwd4jurE+z6LA3x4/G1zs
4evl/LRkE9fj1yM0XTAM3NuszW5Nl1KmFidiKScB7pO6v4nmNCBo8aowz3r4ZX5qnm6KY2Y5XaDd
MjeBnaHSWYPoNRPMD/4gRX/p9IcQ6aJC+mbgcFJxo7jz27GE0wcGZ2hUlGgokGv8dk9fYdfg9QE5
1wRQ9dsa1QIXiKlidmuCQxODj1BWJ4C0r/T75Ba2uvAvALj/REvoZN0g5OCsSj6QJDFqxm4aRPfp
zZboYX+OWusPbfZqj8LXVAtpZZTZxxNyqwWh+iKYMIN6NfN6Au27bqXyim58xgElRPikWS/kHavG
PFBIp/wBLwVHP7qxtc6mQLCXRmi8GJ6YFdVvfvfi+Of5IS8jyFC1g4uAwSfQbhtQjpfu/50qwCXS
a8RV2z8YFvZH/Ss6LsXlEWLmBuf6SrUCdV7DrWJ1cAer8RYM8K3dDBHtVkkDxQZp4zCuV2dzsVsG
vAPPIP2W6kEkrgFOH+e03MePyYtKgh8Yakv/YzJ2YP5KNYkDM945IMiwrxKy2Qq+E2LlVRMdLTq0
/2SDLRklio+LIaxUPjAn4WQufOUuuOGLrCkLfLUhYQykL4+aVwh4glMxb68tuycdaBI2oZ+pRd54
TJfCUUsrXu+Edh13A4kPa0enyCoyXxp9ads27hPfxufAtwtgbHACTcAN0l8UVnldAlkgHQOBN4Zr
wGD4WSvcM/rL9H7fQ8enmrfGNUo+IuWsJn9050/GGPhujetKhmY0H73TnrhJHyozVJHvR6Nqom1i
9mkXsmxdI7VNRC+llmlwVTZGM5rusBTpdEmBSrgHyXSQsfdZVPC1la2fwnx66H6TP7Ewumw3hb+n
y+BzvaVytStbcYHgek0DBgdMwa9PbvcV+fJatOvayNHPuSqI5JbR6tTWzOhNNCsq84zoeDSqFG1G
AdcgNniwieHPqRIApqCqbrMXvKobVm1A5laSlCpSy8Y0aR2edI6OvrKxg14tbmRSdkFt6BxiyhnD
3SGxTaUXD3Hh+KsZ8pNLZQv9MPj5QGkcqwJKdPQn6Psf0a9fI/WTVCzWlYBNsXopBbWR8kfAlfY3
3NE2FVQ2rIKDoEpnChioJrN05vo9t0SjU6OpO9xXBVZ8zjpylN/qefa+pDfu+RKGnBKU+pTjI4WV
6rUQi1GuNsJG9zaF4XXLPgVPPDsf2pOcX/sPMkv2eUd78n+9JT4ldZiLiMmuEsKBPnDTyAumTOGG
4OxHSREhRrCwFBOv8+xRkQ61/xSwpvNnl11eTy8blWSF1xc3rrvCgozqJVfznJG+goTldMZaqWaB
aj6OzzxBWKNhr4gRMk2QFfz+L74M4kHAI3ojEV45KEGRQ9Sv+/jT9GgiLFCMmhHRlN5m8H5k+XjS
r/iB8sBumlzyUzdlcFLGoWZdH1uzU0zMcCb2dTdpjKDIzTgy5ZWIlzWnjKYTTqomWGuvMkdM5NFV
VEsBHV3ANbJT4sNw+Kbwd8nLmUXn5Wj27sh/0f6IR8mhCEmT7x25zoOE2sX1P9HhKguylp0cZ06M
poOUL8oq8jXiiRkFxjcpuM3rcsmgCX0m4d6E5ofRhuMvRpB9R/A16POBniXir21F+oJ2jNQDLVRs
XUQ4gHtgKKJxK/cemZZYt0i5+e7DznjNW/XxcPopbYLVmhUUHZou1CpRKe4EhGgW4EH8nzS/IyOC
jkfxPK2AK0AHuUCUMEwpmmAcMJ9/e3wuy4B26/RHYngBXYarYth73ZpEvCfbRk3YPHvcQ+OLBcB4
9N1Z9R5AoRtWhekHjiunEgiYn0RpZlltRibd+gNt/Qm16BLeM3aS+1F0KHHqFotuFOJRrPaKgjYj
DwDAWk36ufbsbUMp3w109PPNhvjWm4pYCktmFeGAvO8pjoX7IG/RXgenv1GUum61ghDnfWPp5eY8
SZjG2ZfzMiCvAVCY7uEufwOlahhQBLI47/jkqt/frm1RJPq5AUsAqLJ2ZzlsZ34IRL51+Vb6bkoQ
fd4hWkyNpZc2cHNlU+cvsxt2xI+foUc34XZCh7ioVcGJWs3i/4zja1vx205i+KgBIZgmAUC1XG4O
dcODDwCnQjlDPETUVaPm4o0bsn1AU4DUaNCHszhi6c2ktfr2FU+E33GewvaDN1oKg6GS8Lxzj3OL
z2LKgdCjCMFaUW4fGhcO83sk0LVAnHglikDB9VdqOqarN9cDCffrMqKX56N3kpfDk169NCBWuc+6
zMaJTJGU/dGACPjNHveV4YBgbKkvjG6QzBIy9aMutbSsHFd1e8fG9xQxpZn0j1WzFDmtcViGECIv
198dm1PEB+BZM4MiRzSgejxfsPyxgNY4rEwEBmxYfQUvIhgwFrfMljffkMDh+lZ09ouFgyNY+v5m
lgbEz78z05c6gQjhavSjk1fbucrai4gbtYIZmxG0scueTN9JeGGXMDo2rZAtXvT3ZyYzudL1XVZ3
YeWB5kesQf4LbJAzZIamEXeRalymCqwrUMS5KG6EBPwOIJcYIka7OlE+59V8Ke5oQ/mpSMXWM++Z
P9GH/vm7ubCsyYfrZC4jHcInGz7bx3coJKmp3j610y6oCWtU5TmH3F/dKdf+U3IGcVUcM6OHtFzb
mNAAb0PFe88bm95OrhXRwlTOuNk0RazCCoV/UOisU2l+HaXf42A2cMKBwUvSIlYBjyPj4cc10ldY
xVIPUkj6TkIo5Q4ckYcIO+pfHBQtxDY+8nAb9hPCWZLanAkQoHlGdSjWCcPpLxDafhEbwgf5JHoW
1VwITBiGIPei96jNe57wyMRoE6pJrykOjoL/JAR19JLzobYG57Op5ZkWCMK25r/p6UYx4SYaoApl
a/Lp0xNjh8CPssx2X7erPjofYZJQFQBsVhiWpnWOwcG1FoSBh7OKAgyMZ3SHlHg2NMdl/1XpQTR9
qcxVX4s/ZWG4bUbNHVE3ooGAYa+wTuO+rPGgaenZs3xyJIoYWSKPoTJF2sAWx6auLPqK8/tdwlSu
d4Tx/u1v04h6QrAteT3e2DTh+OlvpAPCthY5TOUjN/9usxHa+qduRCzN2ueM3jUVNJXVfYCzqrzB
2cFEQBBhsr/KUrIEb3yWiNQs8nnBrVMiZPTh2gqlJ0TiOCCyXnSaT4Ei1QJDJJYa1ojA3wc9GbmM
JJHgYzEvA2kFqyXp2BpbzvSRuoioux3NKFK1QStWI0u4u6dxCXpTIRZlKqWZHOTZuqfR2HUlxBtw
xm2tlQnUjMW90EKvbFMp5eB2IohN0ZIja+BA1j8ktFblMe+p6igMJmZSEMLD6lv3MMhUhP+2EP2E
4PcWjfOKQdrtTHgLmRUnJWKU73luy3wuxoj4fHlCiXK5Z/GQPOAsJOclWKoVeNP/l8b5OYaUEiBK
bPqjD46HhfS6bmUTgsvynMLbB7knscLFQXA6Aa3hkpgbLUS95XFILM0hsNcwLGgVso17ZnE+V3uV
pWm4yEErHyPxf8f9xEskQSZk+N0W3HRyWgi2bieDfBaN7tNfuVpHTf73WZLQqHU96UDB9boPRKv5
MOPl5e6y66ou/19o16YUGhHhc08E3mthHjesx82XFxRuFgvqfOe4YaLTCf/cndi3Ir48rHM0cC1g
lNUdj2LC2cMvYYhBchywgHltWNDfk/Z0nuEM3PNa/iKZnlmAglfbxGVwMtwThH6Hyho2AAqEMh0g
rurwbvZiAlh4tLfW72LFv1VNhjGumhIZfthpV4Reyhs0rhPisG4fx+kV0OBo+jed74BYIe0DhhLP
StfUlPZ8P3xjuPDU6DyJ1qQfdzX13LS/iuMEXyp/IO2IvLbsTooc229QJsNQFSK+VM5W984SeI7l
9Vq0H2YyG8HgU1OftFCWxJg/IyrGq747GGNnTnPYqHlKKPfTjusKQk+AKgt4iVq7T51V7UCDwHX2
ZTTWhK6W7xJr4w2QtoBp02ajAlEiMs/1IrdUfe3lyqYWKzZPxrB6ixgSdTm/ZPOHBoNTWqQq4kYU
BoXJE+9rPyp7Fv2Td32AS/XrfEJ3Ao+LXkZYKUGpwQiEWcOuMCOKYyg7tejJ1AJWukDfRCuY7Fry
v7jO6BMcfMp4gIo6wokzWHwit5q/yjF7giWftlTVKnuNkzJONsYtirq2Dp82SXqg6qHqTy0TYTVY
oOCK6mmnHpDKUryKAdu9v7um+hOqu0Ed82lM90zjXoNahD/zwCJDgnxv/3YFkMlbNW6u5oAoB0tz
cW6w7oHLAg7IUAixAKVPOeFw02NIhtfeQG2gUaP+r2npP8HNegJGlLECTf6ImD6/s547YrCTMk8p
+AxK5NSMk9cWFaFsDZ6XgNmxB58wz7xAWYS4tIqhwHCphpBYOYRoHpqxAU04tFIj5rRy6dWwbQmh
xVBJBm/TaG/fjXyBM4NbTVm+B9qoKehkNjTYvd1PLQ6BCIY33uOZlVtJdkQn6atAS6eaMsghlKdH
vQtf3HBu1HCdFQjjszkG/wYXM/QYHZTeRkxpmLEjdrCRPrKyMXT6PupjLObD/9wdvlyk5ldAViC7
AVEgGUnTM/jKUyAHE9Z5SUp9gkGHP5LHEgNWNZi7F4mWHPnLT7tVZYOYRclTnf2gFj7nnI+6edqA
iQyCRRRRkEPxUM2M2bxtvcQWd77BuC9mA+foel1HFtGLPI5QdwloDUvgHYfs6OVliTmSWoq0x3Rl
pTX1MJdKCyRZD7MANjBuxDmIQAqfueFTWinJ4z02x6BIySVEZMv9ESOnxXeI2TKJ3cS4cxIeXIcf
EHMLPm6dsC5Fu7wqwBspWn582SVfX/cjF9EYzGswP1WkGIfw2y8W0h5RLaiGdk7v7T22v5cGvhTe
4Q0U45qR9P+j23g0ecmwIeDve1enIL6cYydzR+EfccqXn+hnJZzbLWse5OUOSc2mEe52yOUuRUgc
ItWu4Rh7n4JeE1IEsxZuNiajrXp30JbOGShn/dbDPQGpuIVBDquLJKwl9cpXVazDTZbPGaGTiUJE
ijyeQzwwh1MhzOUHnPx3w/ZL8M11KSiqJWRHrxqZzk2eEGxnBjNDYMthA5PikZzvyYG/tVjculUV
KRYIobVpdJLgzOowL6/NIRFkZHUGc4UvdiMS6/FY7HPKiAWnwPUqHhi2Tj0bulDS6ddbObeMx+0H
vH6WIAO7jY37wkDhkRutORSZVLHHqqZ76HzOCbNQ5hGt/e1aOns0juH7RJ6qrb2vLkEEB04WdGdc
Q/ikY/TUVSPsfz8nG8onxkoaSeLFi1lLi2NOMJ0d6KGb0njgXR4HP00vsDjgVZsq/9A6YxYTNY4f
y7nQrrxwkWusaJUXf+BlXAZsKE8mOpPj4gAD1Z13N7Q4nbAjmyaQ+WqyBJDGEAryKsjLyrLPWiSl
+3C3dsnQ4chr4kSe2iZi5XBZryc7ZYg/zN+SuTVEFDS0VPexrS99U03KI2n+T9P6ZgospwZVkSKR
X0r9v0H3Zb9D7t3NgG7pxOdZlJWe0l8mHvqXjW+6CXwTTu4OaJmq4epnslaFQAxY3URAURKPmlY2
mOtuIsoIJb2a8TyWjA1/xfv2zmdXsBgDr/vOnvVPECejgGQMrINDnc8KTZyaoGSQs13ZQ2KAz/O+
BL1/fmwQLqarIuABfXQb8PyLp9przVexusMKiSRUMs6M4u1AO3iVJIkOa1tyihoOjztxEQd2dIog
YbKth2pm6zrsQ2Pzo2nSnlzkBhpnHdbVJdMC87xki/9ylTrdLb1EbVIBDLcpmopKhCdvWR+B86Y1
bbmjLT67R7t9l1Wz5KWyAs8htTKvVJj0TCfzgNllTk2xu9dUz9LlfM3/WWkfNr3qGMx5budc/+BE
6UQMa+0Nr5TIVlFY70wZKdkKT9H683pe8gm60SchwOMZInQ9Dh+MqUnzjjB2evVDGsWs/zkm7eyu
S6Cl2GhS5aUxt0Cjp5pAQBASrrqEJQ/ykZrldUWFuTwGEgILuLntIHWuESqoqsgo+plhG7R0sUpZ
B+oOyhaUdEKgs581dSfepyWrymQdKdtJr6iyig8QSRQXOjQAicEB8wMfv5T5gUPG7qXeB5UePfa5
37F1rW04CavUpjeE86OKLY9+Iam54/vHsOOEElMEICpJQ97ITFPA/3SSoQAYod+VBIWwG8rbbvgM
zMcC4y3ElvwNr9HVi7N8vpsSgmhdt5h3+ZqHyZS+QwHWmBSIOi7ZDcEpPx02vcnaWpLsVbFhIwwc
U+DtqswLSQNmyiCddk1iMCalVTVQdqLEWth/skDlBrdYvhDRJMdUXC6MATrmTxHDbjj+i/njmbFz
cNx8ZKo22dTEuu3t6wsQBgYmlNvK5WDi9/1rGlokmuYYRPbD4Lr7gXPts8ptHFPmy0008yqWL2lz
AYAyb+D7e9MdjnIBGLVW/GpQb2ZgnOUQFjMUTN+2tVRMglTd/4C14raMNr6yKv9NVVtM8ydnDckF
fFDm+KlDs7NfXVt1YQLLuthNUeTb477R9y7KvdSi7CPIV3AfTnwB56iBQXb3xt77oylxlXxObm2/
0hKmoFg2Em5k+ST/XTGGd1J4EI4PrO7V5QjiC4lPj2iLLdu/OlYZSTSsTIu6cp2gx2X0H2599nqJ
tTWvG1bSrtOUQxb6J/cq1U+9+pNXO2yrzXEBlk6HaQtjt9j0F85BJe6kTey2sVlHH77NCs8IW2KJ
2XKmCaL2H42zVr1H89RQ14KVNkcGWytS7GhZwU7GVIkNAMnJHA4UY+FVtqXGJ+f+B8eCwEW0POkv
xlVd6Ca4OmX6uwkWKPflCykHGS/J1oC9YvQXdWFbA5AREsJw+MmgU8hyiUerCO31dyKaP7cDE1u0
w4xHtpERwzpQjOtdSSwVyas5oeyGx0kCJ8Z9LFmONFyPc183H63/F2+GOnhxQF+gwV/+WdQS6qzx
CKAyZd94P8mPEiJlnn+hKClBERfYeuBJFkDyyGs0gPJ3c+MR2M17U3RqJCb0FqRFj0iKxxMwfKLf
cBIMSmylVnUmRw3HUJVphjsVsRXt5/EubUZ3SzsHLqA0tCGX2Q8bAG8fRvsIKQmva+GxXs5gQBh2
bGpjxOppVyuPaQEdeo72fUZijCX9CwitE2+n2Za3TvyOst55+LxPr6KnQzBNxBplS0ljuKeresDz
3JKUf9cbAtsU1aj5ka7Pc7zUDhHZv8x+bKdkQdLTRONwSXF3JJff+rg+lQ9V5R538IOovSH5nSxC
LiiSMJBFPDNW94dz6HVoNfoHGIpV22blQYxXLkGDdNfCtIziv8bptbDPXB6UaLROd5OoMP0ILoHs
tjnjJ2KsZJuFq4swXdrgBhYqN/xkBlRg7QAy/0da2s/0NlZtPpNf2o6k3Hn8lukQHMpnr7heFZyM
Ud8AdTVrbVXylWSe3zdPZZaL1pJ2KkAiHjyqvUMnrpz6tA/VqW7nz/YILH/LKlI2gFih8z0zhfxw
H/XHLO2EmDC05TNQSL8tptYc/73IB6D2gmmtg7O6GS0nxL3GWJ2GbHiCjByCP070ZirgvbvlqVDE
2u3WwuHJxkyenCn5DPEWanlubF7efog5fDeSe2CWIHjSeYGeXKjSPo+n7WEGvti7lO1oPWfiBeRh
UtAHdmVEK5/sOQu1k29HsdF/Uuo+/cEJ/ZkYNPM1Ks2LAUkh6/ndBMFUqByMUlp1EiCtC2ap2yrX
d87MTVitfieHco+inFOkAAqF8E6zOriVD4As2IXdlldumOiAybp/ao3m7wTnxhB7lBBLxMSpFVoL
72UJgupt1LI0Qm7z9odBdgGz14ni0gLSGFN2QSuGmH7plkmQ605RqziftGdQHFvuAkV0kGNPNJTC
Tt+rD4fSI+UvX3TXDiD3SYgUyLLAuTgxE1IRhkZDn2Q7YpGqsHr2tk/RN5695R3k28kq/dUh2c/p
55qw3MtLWWvWrbK3z/nUT7fah1Eg1qmW1rrteFFeavNtJd+si20sS0IQL50mxg16GzU1kWsZdZCi
YyUHurQW5P55jxLExkzpPqf09DLZAQ6HyDpRXLQ979JArMoBLmtYd3y21FTKBVfcS0FcG0LgK3W+
vrpYae17TVHT7Xbl7nmAuCntyqH+rYnC9cekGMf2yt2B7qBBAv1g35M2oZptQDwK6uDfSRUFDDcQ
nc1Zt2Dq/AcCvuPC6v+krgIvQOSUsP7wke5RWDHgMkx/PMKb/zjxP8GG65n7bdQ4v92ysYVA7Bod
QsPSfW6SAVjibeyWp3Wt3kKwV6Z31gU8rPDM36RVS8GE/F2KntATVyK3+HlZ0Qs8okAZEMliHFhv
WlxvmLlQ8QUvZwysyiXFjGBSN92WSVYXu7CLt+zoJIlR/2p8omEXNXPLYbHKZxZTEz9mB5iDl9m3
ctSJQ2n2JV7VYkqUzsLPb9hbDKzqL7mVGqU4vwTqxOXFODagEAb27dZzOjLYtcmJQ4AlNMhDyo3F
nj6iagnjsvyBo1danqkvwm2NCaZCbe7+OxnIK0R/uajvnq0YXuKOS7jzELKFiyoP++eqmRLGlRyh
WzucefjA24HfzGDIOFcKMINK4ZiwVrmszsuEViHREiB0XvpSzlVA2DfpFBVoNuaQiP0Fv6OaQjxY
coUkH2i9QhAz6rfpIi+NoCyhoCOPaAHMF+4lo42lLwHclIwERacHaePjp13EDt+TU2tRMviuTL+6
dGPjUvmrMNFPNWcn/1Jq8NquC4KIgwqWM8LadkNLyaH18W/yXd7kOaR5X3s47pWHvGURUCcjQX9P
gnKDTzU63rPLEO3oW67LCT6tYc+0+nDwGkzB2LpR2kvlV/VSRWW4CPTG2yOJoIv17b/rkKjvX5Hc
BJOQ9yrPyJTHKFHVWUHNb1Emh/fzyzxwITFGKAgJN/WWLYmW3Ye3bMJFsIYjvHq57OvPPBmGbuRt
wZWFv9z4rzVsSvr8ZK0zp51SJlHpQRO2CydnHvg+2pEjdXx4j6goQWSbHWjD6d3EiiWZylsuP2Iv
NXHje3EP8VBvM5gATjnIretI1PeghhLJ9rno2IrDmrzoPo9X7JL6NStZI7zD02TvpEsn+scKK+Mm
K4KL0SgjAPl/j0A8kEXSV9smk/en9MoVLQM19ndI5IKJSMNZZoyAC9GAe/+kOdKVjuYkp6atsFC6
Rti7APV4U5OwB6LIEuwRivhOp4KRgWCCqF9aXo6MLzhEhMVEcdJ2AwCMr5x4mLp39A5HRgyO4JiF
WwKfp9/FWfHZdf0yVa9nhonqHSq1srKGj6XXLpv9M8j9KzN0QpTKPshxHid89EWrc91uO6BpbaqD
wizy0BLmFM37Tlj9oLGZfr9DWrJakKv4sMlgPxUxV6dLUQsMNc/NX01HGc5m1E/8/ZEudh6JrTLf
KrvNidIieTKPMgayhgWG2aF1oIqGd9cDoVpdfkL4saHxKr2wwIoL6My/FHmkce72KOu7TLn6JUob
Yx5ERKZBqXwLraZ7lzmE4ULuJuXZCMFVE/9todsfpU1RR2IppE5Kad2vEfVGabLtB7sE27CCpa4L
5gXtgMPJcVHEtwUUtwIlN9zCoHHR3ty2xdA6GDgYmr7xRixJIp+TqI1JWjRqv2nARddB/wwM08ph
idzbgOlpRlY0WkJbbb0k/GJ5vO13jKddWBPevS0j6PhVkqu41Z39dc/XDbZjvKRLSiKOeV3Ji/DM
591F/ZCleesNymrcukrVv7L2Q2dZ7eAjYwBT4dQEwmNlud8Pqf4aL9XqlDoXS2Gejqa3DE/cCl6P
XnJ0IeT2ehtE/cjYRsOR89sVJmmPEiOdEV1HUvQgO4e8eibeQmwwLVCzmm6gFonGHGhG/4Fwv5y9
z7+MUc1DNvC6SDhWq7eHGmh7mKykOt4blueb7Z6dpuRsvJBGE7UfJNMdXw9VRFspfY86436L9Mgt
I1hChqRzY9BhHxDRCqIQLiUdrd0tOKyjAoldDwinUxxggB9GKEZ/AJHHUkmsKOGZZWYNK3vbJaK7
AUlzg0PsJihoaPlSz1k2JBXDPq1LNwNn4mF5kZFRi3U7BgE7FZmVOWfJ5tSqDEkiRAo0PWp6Uqhc
l12PvrMatbUplbtAY887wreK/E1mcurboDWiwQzHZdSSUjp5e7OUIjhPSKv3A97WWjTPjRGB/ZQZ
zydMpST0N9mNutMB0MSpFsa3C7Txl0EO6TexaLJGC7C+wQEX9iiVXGiJyb9up6OKtaWEB187sou4
x7yl1Ik+fSA+PASMqR/TFhj34QL6qN6FUZUL7ginOIGsyFWgObh921CA8Hatl8K6mhiiCCE+DWZ5
WgSsy+WDjNEiBLwGcSl/2XS0lBm6Jrwe6lvi2JhqyVIXxBwK9BlEYw6StgXsFdshsXTiRVcH8eXB
LrQ+r7kEZ9tOSreJJui10DQqgYWQTznu7NzhdPolvCTOJcWO0smqk4KgXapAmeCDe5tRPtFBuQX5
c3N9s7sMju7eXy/TSGMXPNVw/3uX9LNH0CzdUFyjueim12k/BcE7FJfSPsOo78YM63lHwpW8VOTx
Bw2V/GyD+cJZtrTXrPH7wUPDWaP+z9o4JI+CZ+Icbb8r6gw34n2yQKYgVoZy03SOtE9EzevLJmI0
A8E+6kh0Yc2B9Co2r6NJkUAapI48CC/HC1fZgZzoOO7GXWK6aJrRr+1z3ngpXpw8BUyjBnAahrBh
YVKHfVwC2zF3Ta21Y/vOOUpJWszXekWF38KB3mnW3cAH5Z1DuM2EkKbQR//kl2AWC4HCb/TIMpck
IVkrRozeIB4YyOiffiE0UIFLalMlewJ8QdWlyIXr/nAXwLs/9H++sNoAoAYtK5RHWnnWIxXN9UtC
J+CIx2tOJIstOseMVwA1bGSnxoymrqrXf0JWRD+etvCxBHkpf9YJ9S47q2HrTW/eW0rQyDPVUJck
YTwNhwKJl1lr4nRbLW1Xapcl/W5w3p/reW5lvU9BLVfViAiijX9HXxMMGmLV2NBFTRQCHp2d2EFV
LLuS9WVdtWpwgmc4O8hOzcHsbCejEke5bjKLaMp5ZyEE41TfIPXyzbp3B3rzimFZu8qIBEGNFnMM
hPYJF2StEG2Zi4BBR4UkFCdDVQobJfsZOhkJ7wzz4zuXxmSWXDA1OT4fOZ0IA097Dv6T2OGUzUZy
DLmCQUkGdmZ9XHBVyEF6drWPfLFGIPmyuVZPWG+uCtiFBgK824+bfQxP6DUf0OVeyAumvFy7rcsE
oe63/Oztx3h9WlT26yskAuclEyc+pk4Ib9CQTY7TwP1tKCBsn/GsbIo/HznRaSSzBpMvodzozmxE
jkwql4vjKdNvAylAnTsVxWgnF4RjgYbzFj/fkkPC++6FoVz6dllXyl9i3Ku0cp6vyJqiPCY0l2fo
3C4I2XoRf+TsVENznBKm3HCHS0Jfbx7qnmTMnE2ndOWWyH0H6PvzaxKWApDTWGfzGRsB8Hta7fFE
DJ0osHFaNwPCFG28XS8F7K1wfelLGlcmLVyzLVEWVzXYD+1y+VGNIi/SChqop1E05Qm1xO08MmBG
YlkbrUcab3feDL2Cir6S0MkbDhJ0kWDyZqCTST35iClyxvfGppHvEBTbNFOyJGx4kmlMGOgufoQp
612VHf/giz11WMX1OwNMlklZpjRMl6l3+gzUjiXRLm91ysfleYmBSYvQFlz9oDup1Hwy19naIUxN
XberQyy1iofGGs7UM1zHo414BHAXhfvo0dKsJvOayKK6DAaQV+QFRFNTHRBet1zw6RsCOguPU0dc
YFp5XJTxOVsVlzunW9COwU3LO7fpvqMJ0w1LC7FDXs9nM3DykvKTtov3TusVvZMuzNBHiB0sGPI9
1FwQeUa2vagralDfacWJDAA4BUzimTL+XknWwzlGjmA5o1nnGCy+HO+A2ovJCVMC7vzrCPOcjVgP
xTHPR2NceyOmsgxQOxH0k0YH2o762d6+rP9+JGTepsxjx7c/Rk142NZeNPEPRzeEaRa//3fA4s9h
qaafTNRm+VvlwI2LJnkS43mS5GP0L8wB7iqZuHDBhFqScI+kLHl5iHZPSkR6TQWNgKsi6Br39A4x
Pzc9MQPRQcjZKBXUcfqflqERChkSNoXOc3mOeRCWEONI1BmFee5h/40HG2TUsekTBDyibmLQSYJM
S5IbHFNGk/HZb8i/aPFmwIMwTVXN8u2Qst5vDYg6kNuvbse0bRMJLE5+V1Ss0628v1cF93PHLtsB
rbtRp1E6SiJieG65aTcl9sPDLDzn4W6nnT3ot9bAThLQcjyAUyCvtcu3p5L1qsOkKmIwuU/a3lnk
tX/YHXU9jdGZkcKe9DQP7+SEsT1bw1MPm0/8UznkQwe/7eHqK3hnBsCCe7eB3M+MOy5EskhmyP7/
zsmQNQGVydk/Fk6/Ex+JZDDBedoa6SR03HuMZS8At9QdEw9cXJDFDhOfnRENLQgjwUPv2UCfbjuc
y5juhmEPh0pMK/ZTAWvi2l9TiCfvytipFCenuuKQhAF/a6V7/8cz8EHFmT6q0wBHWSd3g0viFDX7
FM1UnFKlT0xne6tAhgT1WiCmLSYW6TVqobXulXFOqvgHPZhRudcqvRkY0hCs/SLsd1p/bIyInpL2
XhU4lD7Xk3HhyZxZs7fXMceROGZVMzvUlyt73jMEaGpA8Nt9C0/hZE2DphnWSbhT3WloCSMMaHpW
WiVE7VOnn32pAYMBVzfMOqjFrbKRMHwIvUcZl6PDldikYahZpodUQk0NcQykVZkzkYh7TzS4mp5L
h5CrHpRrnrtq04KGifyls5pzy/0bKkLgdQe1hwL6YayXJNG2d/8K2CCTmS5qUZUQSeQlv2NVK84x
nlTc3qeLBhtGWE72mzogJcGmi/vwMUBrTl2g1L/belVFe1/TrPVdKcaJgiL3F/5iqoLHom6/iYGw
8/1met7tuLR7QMc79WLYzHeO7/zQB+ug5uHD3wVgm/MYZ8qvYakb1DxyjiF69Sz7cH6Q0RhGLbnu
oXXL9A+KGlR04JilGjsrLtjVKx/j0BAnJK5WxxEfG6JgsrtrE9vBjD0wLkyMNoj454hUQqmHAfOi
if+6J9/+cUhn/Y+z1GQuKpn0wJg22xZ1romdojw/fuaJ8SHJ/l/SZvuap/KAicN09LVaPnidL0FJ
CU/BvK10C+ex+YC8EgyQnWU/PpxFHioecqGE2vrprAReQoUdH9PIClt3vv/WbUr8fslH/ugEqCsk
shE9K/YrpXTxAUptAVxUCqX6+Zt9fegxndS5+KzjO+ad2IQrghXg/jmpmz2uvV+i1UgaSM0BIHXl
7yUDZTFz2Q0EuxIA1X3bLfvHDOik++6frMR+dYrcqhoajyK2oDn7LX66B3W6/sUcvSws3NQTU328
bRQyW5SkoDZ66fw0hIflImgY5eoK+mpGuGjX6qWJBzjLg2ApxjGFXWoEKrIzg5ROxUrj6fIVg9+J
PxoTtDUa/NnN5o7XWxn8ZAFD9HYzhw6kcYDNCzcdlPGt/HJPl+H9kSiJCf2hxYh00Sr2tokyKbHa
GPUHMgCbvA8VdLp3KYTJTjMKIaB+gTPQhMpkXll5SqfqOX9g6xLdHYscmaLsnAOmNQo2Hx6wd/66
tCg2RA+C6ahyqMwI8Sm4uMEYuDYueLEG7HPPpxa+dsu1a9ucqw2qw4wStLU6aw4ZQoHZsyYITder
hm2mHetwIhGS+v7cVJYdEkCJHEOVQ2GN6Ry1P3f2+89BIxyRgDEGmY5AIc2Gt1MIvP1PjD8Y4/HV
xM4F93Kku0ZO9Z92NutHGTEWVLdGfbgcOAEq02mV95o/cpGiflDlv+ObVQJmgrThV3QkuaGWCzVV
s2lUmIN53Cp19f3fdtBRMQq3d+ojcY5pU1H2rPLabbApxVFUgK0THIVfb51/Dde7rj1GZVCQy98v
GExoZJJFANr+eSnzR7caVM2REL/5LSZfzGKwyThLGctd7Ve10Fi1iokIVS876y89IKbcZWDwdOpw
J8kXYTK6SwjoO89gXeuJ91ef5G7BCcsAbdoeVTSjiKahcpj6f5RqhiRCpbD/+aFu7x+A3jozebKb
L/KoWGrMk/EOJvyLQOgcIECN13uxjUw2yplu3xF27gKMx77Cvg+ZlHqLfqhSIazP76tQtiAI6iY1
XAFlW81ElMeufvJsTL9CIWCUuDd6YH5dnStr9j0q9XuPiZORgydt/dALtX4FXgU7DVhtL0uhFPSR
YoSLrkOW43b6GeAMChGd3uQ4M/IjwPW+Nu5sef2y4lNts6B5Fbj//p7ymHr+HWHQhZfaRYfIsfBd
v0QEmRhB4/8E8Jn61Bk9YQmeY5ZRByubW169NB3kdHYMdp69DUbAy2XYb3xRM2qrSG8RYhWpZi0j
szirdmp9SXVjIMlgVHHg2MAQv/robk6X7RUExkmSmfMGo0BynNbxBK7mk1Cv95uwvhnkMzE6vQYo
vC6KExCb4X363c5b4vjj9dvePmAgMbIRWetbZQWJyNPatLH503kXek+saS8oSYwqHA6jMahX5Orw
5omJbPLfdXZZt+316/wYW2tNwgbElqkr79/gyQfOUz3f8lDiCCa5jAbdjqPHgyL94Cq+FC+dfzTV
rzfW9B5pVGiAYMBsu7CQrjzIRcvSFJ0xtyppPnD+16HGsE5pWWdrAtYwUt5Qstz6TmTdio4/9vXo
s7OrQLWRpF3t/fHjPkMf7bEKBvszx8e+mZ/MQLmMahIBBgB/rlPs8PTd9aZ0g2oBtA6ioA/+cUZQ
5QLCbtQXhK5yl1qPLqTOqWCZ/MlVIng/eeLy1M91EuMGo4bu6wURPEGymQmiNnxj7p50f5FVIq9/
DLWnIroADXDWS9iie7MgKDn0iBS67GJc8bRPtBlkD1j84j6zEgDplHF3pyxyJfXK9DJKF+k72BHV
dg2VE/9cKRLDtejJd6tGwDwSh9SaMhYa9FfpCDioRxWHCIcv9B1yISOrSVR0CmOjgQVC9QqQiZL+
Eeni7OhU6Y0CvHQpjdUd3151ijK/jy8bZx5MzYdp4D7WKBbItEAIr+N1aysi3kxrjDydTdBmcGTh
4URpMhHideQE6427/LqAMubCY4BIeK9jnKMqdpAOVr/8UQQUcQR6OIP21euW3E4+ms7fwgAmURh/
s2Muiks/tw8EhkCkLV8X8b5OMVk1E1qL4In/Z+flWkxL2n4T36brBCwb0w/r5B2rpIamXif7rDJB
ZDOWLw6et5ygW4rbvqiWT0eXDOILvdaBFMRdnSME8JousVUF+dM8IPapA0EGRybb73IobaHbvEPU
/fL76wxBOaC55VWtl7ToCcofY1Tk/DVusv4PZqI2srTKLIxGk//8V22ffHzhuG0NrGg3tfd2PcTa
HTElw8RFLRuI/kCEOltqzbIdSNQKmPJrHd2k0re9DEtmfvOVoZh1Gc5+jbrzQyNNe86m55RL/UwV
EUYJ2jcw/csq2N29/zoQ4Dki0BzULXPFI4zFnibAtk/u7x695QYhFmLeipHLjRhOiwiJDxv72hlk
as7gHVpvkhJIfJNHQ7PcCvhGmhvWSY0bEuuRkY0U0mkAvs53Xr7KZ/UB6gYDsFTMNOSJZUkkD0U4
sqy7iQ/I4XBN4D9w0AAtKmZOgJyaCC9wd1lLqn5a+Yrwhh37QdeSRr5O3wzG20Rs9AWVbTdeBfTC
jU7Mn4QhhKlEyhDLxKvE9kpg9U5m9Gpi/57h4qBK5LSkzQKAoQnkm4+W9YyRrY1cgdvatzJCfbyn
rtGJKUC6LR3w0n1zlWEvDt1pEGFZDGXv7rfkwCDyTJgiRDEYqWq0jh46j+s+mUqRYmYFNRufWDAF
GLsP8eZjj7s54ZSBLFiNpLtjlkNy0zGCkct1ewGR9/VM7ofcJE2qp91qGwaSRBCYZ/a6yY/Q1Fs5
FA/LmORyLA4FIa6YN9UtWNCKTimhoaIW2mZ0U2iY6MPSzXa2aOAhqHsU2x1DEY5ToELz1PukNora
NNANzn8DZWsfwIoy4fLGmpHs9zcBULM+GN0GXSRT/BApX4VpylKtwRiXHUjfZoU+wZdvRNYDxdSg
p0WoKZKf6cd/XzcMXC/w7AEycjd0P3SnXRBTZW6UXlDaYqHlx5EJYDq9v0rCSRELUhyEXXysfXfN
R198Ar9Iieqc24s+6TPVCRcEc7w3/4U2bYfFtqRmi+Uv8x373QPR+FK9tO7MrK+JyWntlHi/5Vr2
FWV6rNEDOb7w4bhYmxNnOLSC5NGKzLYvbhelMCGrhPHSy4yLxKIPjagOU1chM/hJLur2boqS3X2r
iacGQPEluuNsxnWuuJzLkiOJEWgJlLayqw5P7ly9oFUsjuZCtdoqnhzezq36GRLe85j8VXpGxlVR
gXxQRQGyvS5L2iTrTeQP0VDN2BGigMZ4OOO1rpDSbAtfEfzTqHC6dXy2wpam0CtFKv70d07OHuxP
a5QO6V4Zsf1jUhHV2c4NTLr7IWNPxlBYHrQmPXfzyQ4bpiRrSMWfSWu1MpySZtW3R91hI2KsBtiC
fGV7IbAb1qNg8xdiQJh9/mPJp745yRwVfqf8C6EjyeRpIZSHcJWrQPpdMgypohbyChyc/rc5t562
KVgZ7sfE3j3xE94Ywi3o7vd3M5eWH19rkRuonKiHHk0hMcZ3VozrwsD2p9liqQtCju1mcGQX8vy7
g7jaFweb7ilKhL3PHNK/OnYR/VKbU3TXuQm40Ty8tcQNk1/kWoZ07zfvNegqIjDv4FkqKTkfBCWx
xEriDHYELzj1WJivF2ICGYUnGaWAcG1gH4c+woTkNaz+9Wg2R2wZej79ShQXewhmLLu/iVo5FuLZ
g5ovxL0IRlWg1UqwABMmF+GxhMWD6zPkEAuX5cifHU2Z4R8FD47ERQaq94kgvFM5lQBaCpkSnubf
a170i5P5QrYVuurqK4yEJuXgQcvxXnixQbUsabVxRBJ6klJax5mkswOAVhUcDiBOnyOIj83KxADj
9S0w2lraK8XQ6LANnV+f8l/3QDM6oqYUqgnJ8OY/bnElR+s1EUctXkdww2hxYBvW3LN/+kFmMkyE
CRoLzxlZeODX+l6C3ueagnObW80j1sjyevyhzv9YNQth8CPJ6B9t+EewuHzuG5bZRRi//jP4e+ED
QmvEHuu0CtkN6sKiLKEq9ySd8Z3bKeI3r3q3oSdfGvBsthDoiq6Gvv02KXN7Rkm0OYZoYYj5Duju
Um5N1jNK72Rdg5zPozaTum3yKwZ5PkffPt5aiTKT93GpmjFu+KOGSM8ojcCaF8u/eqH8OlvpQjLw
SNflm7BbK0Hf3rM4SxBo5ad4nqu76tv0Z4h2qiz3RwD+X7S6OJZfEWT6k5XdihsyHcvbeMHMgmRx
MmTYGQ3OefvcHoH7Chk5zh0PlLHYXyo3XLFMH6zSruxDQ/HHtB1l+9RkUJHtuIz4+iXR1PX6DbV1
WNEy5QZw1Du1edqOaX/oQXcWc6ouWXu8pZ/zEoMpMHK+5WYN7dLv/lFDwgCjV3H2UPHDGlFu5PGz
in5P9wOTb7Lg2IlovTFnVYBlWiS4JO78NQDH+6ldOb3sJx4bU+9gEs2XzpEyEz0fnRbxHXabG4rh
6/vuNCMe3/3AaGttQAstHl7EVrdwq12VLurhCpPO8MWGTrBZRoeYIaR0ietGRsp/SrLlRmCR82CE
3EroGQPi1hc61w/alHl1I85yH2UVJbaqzwgDeU2Cd8h3jZdACgwcIf2EaebCjVKz5UqT9gBvQY5j
fWWpcJfU9c8MUhqpx9xcLeXrqO6oUHqTmT6mjNoQKZwc487gtiJUhLsx8lizaUnyL4sOU5oTc7wV
OVsy09PQEPnd1Os2rCUQRJyMrVxIN9Dk3ztZZkVX8xhB5sxyIfPiuTQCa2KYpKuExF5vpm2/aUYy
q0wsziPe+X/5P4xn0XYZ7smnXNIQy840Dxl82RN6o/fLUXJig6Rg5/nrq6+lyPsOrULRvh7cqGt2
yiBs4Qo8zt7BSnC0mMt9FlQDDF+yoo0y0bgWVb+8e2xR4XNyfIbyUZnUKuCeWvSFNakWfeETeHWW
15pyN1z5Ytu6E1aSmhEnlKG4gY0Y5f/OpTrzI6pxe7YRy0ZtvOOaRjERNn9cRDEG/B32dkm/6XqI
DIETrIO6WB93OlD8XF14Qa437P3n7Hh4R70XWla5vwxiUF9+4px3LMoOq9xg/5pxIV7Yw6oCUtyr
wah1H10zYzHJieVuS3TS1PfHCtxW10zwBRR1SxJPcfC/vXetUUA0JvdD9F0poSQ1yd48gqGxjmlB
ZqeGdnQg+zBAmfLWdIFACHzUwhaZTyNX/do93NiWTEJE211aKIRZnKWWrnwdjNiRuyTkIExetfXs
KKXTzXmGltprAE1n2z/gpAzxu+0LL7aPX+i0vD2hBZi2yt21YOciZ4Ccz1m/heoVHW07iS08cdjt
PusJXREhnsg5TsatIVwP7kfTrRIF5Xeu9PwjmCusYAh4nOXEH5jYzRXGMs1IwvF6q1GeunqSYcip
Yy2qiBiVKzwmAwGJJ0NbRwq8jGYjUR1ddw5OngE6IhHDKLw2ok4rXK1ydF4jEf+YyGgDDu9QaxmP
Y3G5/NrSc+/oy2126YNON3DrhMEqLXHAjwwA2l4odL3BFujG/A49IWLFhWPaTdnNdBWHp+RlqQ59
G2JOxX1yeJEYLfUrRpgBrU/EaRwlPPdL3nOYzC23mTNA8ZQeE5vSSmC4yWfITVmHozhZifw0FdI2
YeTSCIZ41PbcSG7N8/jjArOGj1wqq3MvQl22oyOzBLu8bVrch51QNUZGxAzNWuOsPZ4ossY0gkTh
wuwaHTtbSX3PQrij0LWs7YjA0unAVxJlkG5mhikodfhD1+XDG9g64wGxKXpo/+Z++AuBBr1etElZ
6rHo2sl0CSIn9NII87V6I2gTCdrmrOXGJa+EPILa7HGAHOWM+r0hm5Nt4vebllTxg6toUn94eslu
GVUW6B5KBVR4RCybOw8eTDXkoHg6MWpyLAWdZoW/I8Xgma9y65Or7JyM9Z7WNoznvCjOZ8WrF1MB
Q+CaowJeWKFWuTimUYrYiG22il+CK/9wuHmT37JKbnXvQPTI9bnBQKIoCRH5OFWBiYzYLLbjpN4L
OzTG5qovKAg2Vl0NkJmbWIhFyG0Gf7PBbFsNX6vX+gw0of6V2rnYHQpSqux1wSFNjgB9bKqwOGOE
Rr0OaBT+nIQJZVr/7o0vs/Rlrt4GI0rrwIS44s0sYsKxDDFrqx5r5JfvcdC0pHw2vlkDfWXVxfC6
2/Jp1yXSwqu9zKsGJBoMbpi96SNiohFjq5d0+I+6dfv5e55ESBk1YuX1fUu0YscVzr7hYS2jrq8F
7jzGRJ7ovEG8VCqNLU3B5rXzssKJJBCMPZLlisJGkdAwvwAG6Ibzg8JdgjLGQUtDKTXb2J0Du/ZT
WDuo8a2yd9SoQnLpPinq8f9J68EY6Va+oiiKxEpr8Mmby6diQl2nrFC8I8DQbPJ7cJpZXzZSnhO4
f5nQC24pod/EpWaRbxP5+G6hKWlVEifc7S2YQNnxVOAOZhOq/E0LdqjBrp/cT1pWyag4Fr0gPNBe
r9CUchm/Ilv1NY8uKWtoUg5YK9HAoju8pizUgDmyxJlmrAWRzHuI7y9h2Za5ssWdLZ3di5boHOxQ
SXNSs5ljhRL3S5JuJuyBmw0ve+InZGsJaN+99+aUZ5ePTjgoy4gYZEzbNSIXWmSSGLJmPghda1bq
tftihRSap4ePBv6gkZZF5lW32Ex11MAhZWcr1vpjkg6JMxxnVVLKz58iBl4Yf4Mkn2oToS/GFAIY
V6JiClTpAexkknqvteQFbOhdssuQ2TzNdLWrOZaAFakaNaAruPmsn/TElBWAYdiX7s6P0uFgiJlx
OP28Y7FwHUoPYH0WQEEVFxkvnsUWPjzodyIqzXzoG5pBdLZTLgVkxZnNYpT1JiRNEBDW4Prt69Q3
xIPbe3mWBp5qrKd2AROe3HdMw6PMR+FbpGiHXBFtgy2203SL6FKmvc1oAHCXaVOxnSRf/E5/OJxw
m9o7Domrlus20+n0hMWJn7aYGexn5rs5e5yq7wKmFe/L1Chx4FtaL6NQM6437QBKYcFWTcpbpX3U
BJIQEgijK0eiFqV2qp0tNW9q8ncII52jOvGMPyeVFe2OCzak49BNIRjFwQuREwwsHt7R4cPdrplM
s8L2nbGwSdBoZgVUwIVL+B32EOkO3VhuLa+hLMvkuqVKGKKDAvagJ0sf/yBSDU7b4YQVNh5/uqpH
+AHGzx0tf8AU+jFYYHzITdrUnZTpIRbY6y3iHZIvbeH06H8JbRkRskNcbhxmW1QNZah6NLPG0IGY
JLsBiG9/rg1PYs+FSjEUknsfjb8LVqd5Oz0MCnB0xCiKxKvTlR8CLMFRz1ptBtXlGnuqcgw4U7Vf
S/21bknAEkhOUR5ZLE1MYk8aQ3viLx7snPvvXNq7hJYuKAi1gAadk3IvoWODPUBg2/FapnqMW9Im
LLESSA17+ExXmqzSHXfh1+SKLNNKkt6UGEFM/kgDixxHhTefkI+oATzVf9t39Bbez/ssWgojPR9e
SQbzXkGgBigGb66FDTMpkAwReGoxwGk8upkBdJQ9fXJ9CnHr4Ri1eRWj+b2rh1BjCcwrhQkKE+VV
eZXF1oQ84zifVQVp9RY/EfIbPIvcrQa4wR4hRD79x6nY11hgglJ1etepO+vcSkxGDvzy2vP1F/1l
j3YXxSCiG72wmPpWnvb5fKb+gpDHEwdBCu3Yl7tcdru2p2us/7iqDlNK2U7uXqrxhrpHh7MpSR7o
vO94OaKP0FrhaU9XJglA23YOmRnoaKaT88YH0Jpdf5c90RXSqawy58AolUpWk9X4Y/FqQczl61Km
Ln9Ddgx0a2pitJUljcwcBjAoKm4+tmxqPChAfLIiKR4EZVf9jjqbpO/yhI8PuU1gVMoELpjo6aQJ
+AymDASUiL8kAWTlOcq6crB4gmArSNKnoN98n6gLwaejL3xy9q3AeL4vVp9HMAymGoJ57I3dCRpr
a3HFoQ8HQSvp6XL+4RvW67OyySKeReiL+bb+gd/2/2GwmClbhG81FydnSS1t3C1LrZbMXYX72kxF
eXBcSVSsFbo17m7Fu/AcPEEqFSCQ2GUEhLBeliDJPkeHMRibxcM7msvPK8NlenLSRPYEQWKf/+v0
1B8K6Z90QYFe9b/eg5Odm7zDngLLWWRvNc7np467i0jGqQNVy1Om48DQzEjcZFiI937fVce3dnmW
6Cn3jplOGeHSVDAhsu8hgJSJLPGUkwaYli3nquNb3JHXyiajhQBobT4mrjqW/aJJp4lUyrZaBuFk
/djOZbJaBmKuAcI9ebqqUTDqJcJXt/yOxsLzK3kAwUcQm2xUw4uw9jZw/PePi9+BtStL+Xzt2ygQ
0Rej3DDEldnTJtJ2O6P8MDv13CPEBNMFIrj8PVGhV2+LxJJ05y7WfJxMgc2Pnvq/fpizMUCGRwY1
b42Yfgfq2XCP0Ta/uXtmcC5+csoxUhT0Sai7BTQHxEV0VkN40RwbAXAX63wKksULIaZ36tswH5CA
z3nDm+Tn1iQWUKcQo+MKbXNoaBjLZDGXUptYfevA8gPpI2GOeoUfdR9PPOqM0v0gOHfIi2EKXvOv
sIWtDlzUt1IBtDDP3p+I2WPPUH3FTskI1DfKBhYA+CaXNvWJBsIChg40M9JMH5YONlMWgMnLA0W/
AuJfYaHukFZCbcgSzzQtINM1Oc9ygpTRWJZUsrt6otc4f6M2GcZbDd3l+TZtpQ0ShuxweA/7ZLpe
1Cg+g3B2nIs9WFM1SVpSp9f/jLKn2mGMIK0WSvI1zm291SmCDSu69V0xDlSIp6iU6cc4QLa7tC0Q
OdyrO1RDqEAefsxQmEJTjbLP7jo5visCKY4TgmXl3l4rJ7a1pQ1+CeITxuJRfFwbW2WFdv6yh3+T
4Vuz4BmrzR4v26YFl7vqv3fBBtwhSvJCIsYIFVYZCzAAuglMxx8W0+2d3QvoMnPG2KohircVl8Pj
XqmxuiquRQvFfz46Okiwc56Uo7lx4JbfHqqCabfkWflGV4NJIQZH97CX/SQuUauwCv4OOPkJYYg7
3bQYmKXxUxuCX1QaY8ecJ00WoqF3fz721oPxhh1Th1xfR+U9b9Day3b5O92hI0l7YXsVAABn8EjS
9dVFqpmmmcdp6nbl3ko19E2l5Iu/3m7rIzWLo5CMM+pHisv4VFXDGDvHj7DIh+M6xzBhdJlrC7bc
7AVFujisfYHT30JplephLQkNvGxBQyzCbvfC8y2oOIZUC7jPVyEt3I5Jav+qkl+CroMfNohyxuhd
69LD2qRiEDaMFaj1TeBXzoMzH/AWhlLrzZdOBEWkazmBwNETCcGnAcOV44bq1yUHC6IIYBfXcld+
8FQCZG65ECwuXVzgHaWnjDQ/PGFC8NLhFnFPl6dLpHMwCUmWCDn8Owk2C2FxNPqFGjBGjf6m5tzS
lyDaipwAHcQY1gs7aKgmIy/ALe4aRZKZL9ux/eNvOQP9ASjoIgSeKMQeaAPlE2+Zo6rPNBIFMzCK
IawW5mA+0CvK1eH48aNiJxKt1g+w4iYKoUABDEhQB+/vHK4C5qunfkPbM7E0rRDKcLeF1YVjmYwm
MLL4Y4TmizC4N02n+W6VP4mWRnCHheQOOrmixnAa06J+d3nBm3E7jNZXoTimpvJ3Pn9/ZgIekBnm
ogTZRV8xt4XkYzpEoNeBZFZgVXe3TSBSVJSkLNtHIZh1qxV74AJ/XHOcU8Cxr0l7cLD/U2+Sk36a
ByLQyFBkOHcHa0E6ejAF68h6kk8iORtwJH6ipvYOtPYpHasP36donzaayCkJ0DnQxGV9hZC15Gca
ZoP70VYzHvdigyXlvPDCBy2swLJuQxT5/3W7rOLkAAIlFrL9YE9iap8qvt6gGDhxa7OkUewUSj0q
333P5RymrXAXilaj93OkkSLHARq4CbouBdh2HCr2CA8G6V1lm/zb8LL4rBdlYVYcOTMU4Rj6cpXJ
ZeYvPoeJ/r/01LwHPU7LmNIMEs7FAxYwGgu9TjfpKCJzmGXy4+39FCSj2lkxRUj/kkSrBeBWgg3d
mWHJFFAHUDD+rH43I7nde1+9A20kAsG2eyXvpdaO1bFBCfIyzOQb60yXuVdmnvHHeUte/aToRqlZ
L/DmoRI73NMn7ANNp07aVxPseP1WufCpiIHknjWmWjlCylkUEZPINmVqClFjwxZcwnhXgB89rLAs
ls949DTp+V1z3Fszlp0gjLKfXMeFSU/McL4JZ0b2A7rMKbJsQxZ3sMyjfcWpwk92vBm37z3LbSPV
fcL4yQRTr6FRSPAGIMrvCttD2vbJavLwHyyJlsQAflhRqpOdHIX5Wr5mlv6mwHfk9baaKlH+OXJP
7I0vD4e7RYwx1kQKh/fuIkRtZ8C0Md4ic1p6LexsMRW7o50IlYeCE5Ukb65ejTrQP2WBBgdbfbXO
Lra5knv5K/5YEwdeDBp6a0LX0qi41m27B9Hi6pXFBfvIJYKQvy/akGtyBc9ea9AI1iN2+WYlYfxr
Hbc0I9udy8tzT3EsmoWzU3u2FnUT5oU8gXRwJQQED3lKYu4HrtLjmXEBTNer79zG1Q6rE2UeIjaG
ZG+7LNdSRPujg/Z7JQJD7Pe/2LiAxnefpxieOts+J9WtdPKd8ipS37Z9FxAyDaNMR8SZuSOxIixX
5pkk3CLupKE3h4DGb54rpw4FPmn0PGtzYutoFBgAtJHXQOud6qxqp6KVP7S6v4Bjpd4WaIpQcTYV
pUSfabNnhbK7xs1Cb3pahv/TfL/JQirD4bzsX6PsT20qKZ37I5wpvsX9OWtABfkgPZmG6RrtT1Bg
javPdSs+DheAdL85SKtWyFb5MMyRCd9BxLCmhAOOxf5KXdJZQFXxKdevUQOMuQY8kpS6yxHX7nLp
SWenpH+p/n4LKlrp+ZCJcdz/BSWkYPsp/tESnMTJsmApckx0qJSdyDIJYBjvHEY9OfQpyQCtmOIr
0n6+3p0LRfXw5C6QUeogBYcEworkreO8ER78Y1H5qWWlXIeC3luEO0tuZ36rPggKRp4xbFOFXW9R
0hE6sKHLBSAVQDwWEoJ6rD3V1w+aiMJme8btt4J4/uRmgK8Xz+SPhJBY80XXCmKpRKxI5Xy7l20D
pt2soArBoiJstH+d4M44sXu7cJGPT3UO/w6IqdSzLWrFd5ZIbMOQKOwa2e6SATSujfVGnH6KzB70
zlM5h+34+bCpNAHzTX27iEQS88vVHFEUm0QdecloAlss0ZPFqMhNCMA5meHrul+ep8j+cWWjTMDf
0C9B42G2Nf1fi2zcehc9lJjNcwWu98cfmLkwdvIO68GgZIQswNvVSRQkm5tqiXK3SFXhQZh9lCGR
xQWWFw5cwQ1JTJk0CSOFLeWrqzVGsVvw1tIKvwwJnC1GgkjRA0Qt2IgVwriLHSDSzhgjiFFmc5th
mvN6nSvcr/p3PY3Xh8bVipl5x1//wODElPccTLIWUmiue+S+PTDgCVIFQTRGDDYEAGxh5KDkoUK/
7T1O/vCma9fYvhDp1dnwwQ1M2EMbiG5DjhpZ4GiKLSIoZxsAyFWxH/axdaCYgrXdMBCkzXxu19Ga
rJDp3Ux2G2MSDWOf79RkNJnWrmvYrjWVbKuUE1671P1/H9wUYLa93dPFXUmcyA74e39v+eLWZ5kj
N3O6gF1mAMGxeToHSyL7rUDC6exne+jtDL/okfFEpkm9A1+Ra92wggt4rcsemasFPWL3SVPA4DJA
Q0dht/0Pv0jhDkCaL5QMldAAsnCkSkTfZmz6FsuiFypowJ0jlXLnmPcvrYDFxkFUQGpm3dj0pPWp
wUkfJMfyyABSipexVT85n28S7L0dIxHBoVQcaN309HYvscmTRvsjS3w/VsLgEQwtJMF9qM0t0Pa3
E5eQPNV9YrhDn8B4wp65Rc2zOdJQAAgpU5uMwXJD/OxUXcUDB4WZO3hmtCiWHg0SXDElsoUQT9pS
CEZ2nO4D2M5SJNjeQaZ2uc2GaxTYMDItObiPBODeobIgu0rewghMKgDCLJSnLsJH424x9al5VqE5
Ho8SiIMQD2hS181o1hGP1eUoQtCPSlJl9mUN5ia9vGNAoSygkNyRAm3nrdvy1ae0RfNBjpYTBn0v
D7HkjxgfV4ljfHsAiEXfowGBU3FejVWvgQb+M+HJFFjvkmi7kcd3gWi6wQqsdeKCiA9ysFglwS/e
lm4SmaAhDrcIJOS1cAVcSoGTIXY42wd8Y2v/iX9EaujtBhA7TwUDoBkriEGL0QzJtFZ6HNf3H/35
N+CzjgonJYl36inUlTb+qXwb20uygPhL57jPUG9vPBIi2G6z/G5TngxnT+uuM9reOJ3keqJ3Rieq
Jl9IOXDv2dGKsDyz+McWakb9f817H8sR8igR+yhr9rI+GmUVdgPGhjDi6I0puols4KaGyy7jaOZF
72MKm3hZVwQ0rimLBSm42a1NYj8cc8HBr8DdvgrJNTA9Q/PGdbkS0zlD6Hy/7IC7XHBWdjbdz/vI
EnSW4A+lXR9ksZhICwn7I11CsVrmDhdFdiUmfIBNXNa28oH+I30gP3ncp2BbGWrtfMH/gThjk5wc
r4tiWQDGLJltpb+K3GI5+i0R3SLBBMpuJb67cYqrKfttk0XJOBzfi/jZDSnY1sX9wIw+YwYwUtMG
HUMQ04xjlVp+xzKbyfIDZkyve9Ejcv0L3Fx/EkeWPRWPwFQud95etcyG18j4gpu0uvyunG/qb9tI
XyywR8PzuR6PKDkcDliiTh5h1ZXHiP7XAk3tXqrl1MlYBI9aCMIWc+EBk2+hhtt1f2BpRhuwABTy
sXLMpTav746EkGSoh6I++79xHSCN13C1sJ3WKx5fs2zkIuUKzsQTmrVjqz6dNkqTgfLOuaR71ITL
LQ6c0Q0pCAeq44VYwNmvqFyUfqYewYAltM039YFEsNcZghHJVFrI8WzoFX235aaO7M7RJ3Fpkxc6
fSEO+nAioxJLrR63eWmzrlRujNhobc1Hcaf1+C65j6JYgldEw1I+WFThccQoI34vGps6I1Rf8Cct
BR4aOOrIYb06/gM48prlZr3H1dfm+5S5G1whd0lykq9kStppZMvIFmLDDRB/9QjUIRFuaKuxQiL2
EspE/w49SO6nWh/Bx5jlhyYUfu/+LJHMo+nXYOTMTay8Wg9/dJgu6d3p/TeazTlkkoeMjwkUHoA0
sTtrdaUXz/5HD+EvODucoPwCt460Kl5b2M7MxZvwbjpvcR3GBaznBSzp5+I4G1lkC/L27CIDBbgm
PgjcRdRyBgkVglFH+bA9n8oki99AzpSWNXmIHM/e49cMElgg5ZLSf6gWb/2zahL0RQGSwbuhf2ox
y/T7wmYgX3Ofx1U/4iGAemmiAeumDtBlR/gokcFWMaR1LI3aqf//qQcuNxYp2yNvAD38tlwPhcUb
XiOQv9FearPDqh3bEjfkhN/IHI+ZHpLGlsys9sTX8b/cYnepRKVYejAdHpmnuNj83FGwr2hqalVC
qCI/+HqTCA6HCbcSPlrYtrMtZINeyzbwflhRmKbg0upQkwm0W1ROarNXxVyEzuzG0VQ80QQvCpI7
uZOvRpXJ93o6Rjv+R6HboE7rw3bUp8bvAtbD17IIlwEIq2L5Caj4P0MF/TRArnoF1qxsjMhWhCLw
0VBu2tGMGIYXw4CvAoKtqCEid2zG+uxKe331B7Ik+e7tBqOozmgcS0KbmwD9DXk8+5EnX76wKJXR
+Vbhz6d5wRNqhrcdGxlPn4v4qm5dvNQ/ook4ktZB8NZt6wNFjJNnnpV1uw4AXw8oGa7nqlOjMDhY
r0FlLCLBd+w7ohYUjR/ZMf+33tSbDRO+xF1CWZFCfN/oIgyaResA4ujHCKJXO08ICh7RqG6o+XM4
P4A8cmVHZlqVYWRjCRvx8naxqAaxf+DiAGm/LOUMoXzcprEQ+xeKCnTp81QI9hIxZe4+7gLZXyOq
A5XjUtm575jh5P66LAQKQSsW/QpaAIvj4YH5AiQ/iTzM7SUlaEzT7QOvafpSA0npcQWln9gCQhcK
CR6i4WVklhYfu0/xSQPBYScDz8Mn2JEm9vRFDL0j6Z/WVL6L70dJjyfQx4b091f5lOTsM8FWqTqx
AFKLRieiM18Lw8SDBZpLl495HW5quQSMeCYhtms2zRd3ttKfO3v769GBkZmWvKMQ/R/HVK+FmKyi
155rygv6LxqimTl6DGTQGUwn2vbOej4R224SHamLQ6tozi+NFJtECUAnEMguLwwkswOoacynYJ/k
5fawHZOjgU5LwzfoPfa8vwdcdviE366mzWOXqJEg5n/WYy8K7b8PO70EgS1ZwBaYWYAFEizVBqOZ
2QvuLJzSrQCfZsgCEpthi2PgXB3BhdOxmBcHW/HdhQd0S+pTF9mi78GvA5HHg6kUhXneW7/Oe3bi
ajF0Bv4hQr5yrLXLwxFFS2lb0rT3NICovjdQZvDRExCO+DfZ9WYODFe8k1tKXn7ld33QEyOiwgUl
LL81Yd2Jx3NsJOf77XbwqzRdP1M/0YnLryTQntdzVXH2UQ8S4G22VIDGwcKBGd4f5+TcQhffCr3v
Yumgs+C3psX3f583PTxb+Cb5aG9VtsvKstF1qYeariZBjlLbkuto4AUEJBC710AapVqk60nZN6Vu
QEwwD/TKTtGtZH6kdeAMet3oMt04P9h3C3y/iR8sKtiaD56hxO9/6dbhbYnNp0r7Mp9sk1BT8S42
EvkGadydCPOKsQZgvgurmhFvmnVJKbDihOpUxdEvvo2LK4BYtEeXVxV888E8Px6B60wb12MznePJ
yOEn+sfKYI8Ad8vFTKO+0JL71qSEG0sMHed94idcLgGoJ7UnrlDVWfkCLKdJZBYW+eCbX8tyDk04
It2ZeMBrL9p3qnPxBR7WzwQOHmj9rJmM97p6pT2IT0MJzalIVJoZ7PsQNSa//L323XOlBdPaSLsC
y5bgT55AAGHfQZaZjlMnBinPtL3P0wPwUsffQRNvRXqrP9PnbADYrSq+jxup/YtIY6SG0jHyaWB3
cIVXMZ43j8qpWm+a6Mp0eotKPIK4cY6z08cGfC/QyFFc2q6dkINmVEqfKnjuzGeBK7jluj0otmdU
4PK2ZWDplWauP9YkUbohwanY+KEodoxEsr5wEs1Z7tW7nt83JfSMkenVBqg09YC3d4qrkqQ8mx15
Jtk+nbcaxGAuL41Y4yh3UpNzSijnOIhYzg3nNIn99QORDpuwTHdfHVubfNczlUaqnq8aYT4OIr4K
OthSNQ8zqlKaTaGa4QrpB3vel3msP8M9MWHI8/Ex1OzufNiJCNwa9WpTwUVvD33dFdpDf6AiYYrk
B6cAeQf3GCkiKD7ChyuRegsInOVaB039A2HSRTja+GzgwE+J3lbxfjHG1O4lomlzcRvjotnAm+Hr
+DDN2ErK0fMCyhO8niQZ/MFmBGCUmG+cYy43cE7bUofA0qhWL21J+YLcKhJTtXant5vV4ToOADmS
cfdQJujxJRGi6iu2NGr/2sc3HYOVYuJg1wZZLvFzibN9uPJnlZiQWXX5Wzm6hPY5WcHtXmqnAvqK
yFklUz05aik0uT+9kwD3u8tkJBASiad+e3pIBAd4q01l3Wax5kldd00xpY9Tb5d54/bfN7zJpllU
x84TebIF3e94BXIreR86d0n0oJKz1IV+n4pkpxjtYEMamea1TfgWWo54Bigy1FsTa4e7EhAxuXXk
PVNkTolQ1UBpnwD2Hrt3WIAHg4mkzYYCAr85xaU3ZU5jC2YHz4u/EswRWkuxlttel7bf3iIzAjLE
hSL4WBI1hZPNvVjdqSzUUY+aujF7VI+SHeZ46erivVDekJWCOdDRGKF3WJXvsfMqucyK5PpWEZ6Y
C1vCl/SUIAx8bGYOTDa5EqqHZ5INyZfXC0BIVAF21mtLqVd0Adxfz2sachTTzOO62/1HoEUogfpn
bxQlElXtGTbEOvY4THaXdHQAw+Hw4kBh3MrkvacKx6JmDCaNcLBZMzXM90ZhtmoIHn+G7XxwqKlT
KWBbJj7iOulkQ/ovCB/4w6tPLAKfTq2/kveDFODSCcumQFrRsQ/qc1b1js/ZVpMEFoxHRsap4uSo
oZX4XbUmd90UIoCmy0YEr70faNeFVKbBtbSeMRbOiTOKgB+cv1MHvAFn5CP57QnQn1/ej3eoYpZI
DenN6QfKebvlgcD3m+wYrbixOsHgbzeF5RSLW6oIytjfTZSwjrsl0RiNJlxWCMDc9SPfy2Lo2NOE
Q9Xcx/Kg7L5BZR254CnFp2WbrCmkF170I5UPPIkuAS26PTml0lvewZ6ML9UWU1GZJ3zw8HMC864S
3CFgBUa1w1vaG//lW0ejb0VoKbPJ+Q+ZlIB6sVlvvCf9zSxtUb8zfhPANp3qKwMGi8BV4PrKWJZL
abDRp6vHYUNUV01SVKCXu5dkLCOLZnoHTJqLJB4OPMErnLcewtdSF2Wo5WO9lXyJIXbWEw9H6rZo
S81ob+3ko8CkC2A993SMFqLtjTD3tZyr7j/UrPIqHPZuaDz5HzEqYaQgJBAJueo90uUElXJzUsfl
46Y74Ea7O4+gJaZEeyjW14MYohbxWAULZQWoAVV7XCa7BYe+eFIRZDrYl3ZuLKedlcvweC4R1Eo6
A9v3beOzxahtO3j5JAidSytq9w/ThpFbe+IPtjESLbiZGPMusfUyN1ItKXzCP7lbH4cvOdkrAAJF
AleFU1vgsI/ENo7PIaAeo5osxVO7tSPyjVySL193vVBg4nJjN/3dF8hXx9IUTsMiIPouMXmYku0C
RrI95exKbW3vjHwCEQNAQjikQewvW7L5BAdbIvXk2RLrIiNTUIQuu+xdpb/HZcbZlRIxev/ptDzh
L+TOd5MTyPdnKtUQTTjm5aPRE6kf+3b80cpUm7Aicck6XBWaz4DIoxFY692Iv8E8u7N5n2vqUFXC
qoRjCZEL23qKhjX2pYiMW4L9iCqrqljgH/K5QX2kv7NMhUmMT+il8Lt8LqM136HvEN1K0+Ev7qc6
JdgMERCIkX0+RS0mVKIBTK3O4KhaqNBU+ZiGbmXeF2atWYVm04cbe0dSgBFSnahYghVKusaJ5eou
28vLh7jea4AE6VYgzZQRglRTGaOqJCuFGxg4+fhggxopesD4JiyFaDfI58ncKYtsio4bQarB5yVB
AS/mom6acOTFY8vsic/LykmrbNjG6yTfFTOnj2fKt/ElLyEf0Ss0wlTeaMx378J9iQ+1Wn07gDUF
rLCEKZjhXDYqzpzzSz57dsyVzOaFnjpoWTGgtpCpJDgR8X8M3tHQ4c6q2n7YheMq5p/C7cQl1TXw
tg/iyOdvHH05WJfuNPR7PrkDyn24mR0ljyXEfE063b5y1y1nSj4TBLnbRjtzhzTrnJ0h4awdr7mR
/SSwKIS/PUOEx7dcGIclRHYgqCSWXNRAaGNk/CjzvPI2Dq4MPO7+ad2AROoC5aPNQRN111j5/CWB
S+jOv75hoK9l/Wkp072Il1qU85ire8CTmI8XbQNJ+y0GCtA5UtUeUWrasEOP6Vzm99bi2xhHQj1k
Mfpp9q81aYVCmKYgRAlXgSHH5HokapJdfdhahGIJ77GAMxHj2qs5fNbT4L88rntscWFzGo6LeanZ
OcGTy76H59GGWp4v5kHURPRDGuDBn7xbTv242XdgZrjkDotRWVfVZbXYvpWXPsyRzMHD3smuJOL5
kmVn+sBT+uj0LxRpTKVLzo7+ptL0oKnUbTm4e2MosRFK0CqhFEyPY66a9G2hcNoEXov4eQWMz/C8
wk8v7W9tOlXpltAHV/C5odtWxTKWRmibvRl1q9DcvB0uJAfHP+DLDdK31ME70uUmoLc4vRhYSTwr
duewLXwY58oOWG8cfPqS/JTSuRvCPUARZfG28ZOiYzb8Y9ARSsG+62pG9bBY3aqF1qtI9MigzZQb
Ch6/SyWg8NVSR8h2ndHOUIBNGyHZGUp8eYZnauCZpjvgW6s/7ZitOML3SHlDfPI+FJ1NwCuqKpGf
dgxll4dazEsVE5f3OTxCXDd0e7VYlS3m0L+gRSRxywySSyIIkLsMKCqOLyoJZ0qeT8kuXT6tI46g
B+ggEexHKyoW8pJiniRqWdlIDEV9m9xh4UWXZ+aJnqkj5ySmJISy14QRnFWKR1iPxV6X5pkoIyQ2
RuVnvxw2zty2hLKbXtTMdpVg0cUGMhjcsGebDxIIvozcHNmP010RNUBF6PjoG9TbrJfLaoJ2sRNF
aXlCotbxRlMBb5wEQWuNOeD6nsfHbVgDk/+sgGapIWg1hLfTndZsgraf9p66Beqmk6JVENmMPguw
uiZU9uzf/zHXkBJZyRRVWJBJU1iaPPGCq4UcBQM7lBgLMlwVqjM7dyTnbcYckAxHb020Jz5ua9tZ
rqPwq+33Uh5yZfy1iM5U4vFGN/Sax2Zd0fkiVxwR6TC2xfbChFJhwE03BPZFrTJghyH4rbYQJ1kZ
oIa2ZmoskFbD5G/FTszVXViC+REnzbgaoESs2Jp+lhhs7TEFpXJyV1mu74zbszP9FaOkqQIUdwYz
UzvurUMDlzMkmvTTW0Nbfk31qrVrTIHFWTLflHydaUgUYLU2DUVzR3FJzUoQA0jgZVTbaBxP69MW
Jt/2WzFCmwY6EUfyXdt0ABusuaGc6Dps2SzqAkScZ5BQgO/TBWvd1lRH8lfsEZYsNoNW4SYBUQlS
aKVCi6rFHdiKP6LkqBaNlVmaHpOUkUq19PrG2OSe/vJwsXLJLhNYM18yc5Bg+KAodjbTeK/vgk46
LRgb2oUWiC+79cgFselozejik8MlS42lEU0vMxu4QokooPsJwQiNiT6BbfLeygYqzavccZKfgLX9
jcJ0G0gGVJuh3Qnwuyfiy8zmNPw7XsPjAf6NxqfAqylItRnULkTqV+fT819fQB7oYxHRuObrTOi/
t3prSxcn5B+ZDI/gdfp1CLZFuiPSN2faxiNRkqRkLMi/D4CWYqIMtdgRWTWWYrGdbXryERmMRfs8
eQPp7FteE1Ber3iQYmkxglKVnfw0Wbbw1tMMbw0j+WW1I0HlK5v87ogdqBBzBkqG8AFDMfVNBwJx
w3VXrvP2Y3pQwz+fQ8ZMFHPfW3hoAe97w4J889Ce9BTUenovMxWBBFl3J1HtsfxbPApfZPiEpKHC
LVsbVPNYknLuuMlnv1JoyL9P/LxblXDmOmmQF+As3k9YBBmoLYfFiiJueIVe6pu1egT3vCfoxWGM
IdX/MFwd+DzHea3qZNTE7LszyYiqiia4G3BtFnfnRQ+HjK5sYhhsXjeLa8pVX3JXj1yxRAdrJpj2
/khjGHzz8bxOG5qt8GQXUJbSe96WMHUIXwb5R1mCwlO5AgJdStD7WiG3OIvSgrHnlKspApZMrs5a
g1yTlymV5zTOzii0EPOVSDpPID8NRC/AFGqVfwjmd90TnEeMfTjYctjfkhIlWdQWL4C9XEYnVVKo
KgaX+0hprv+O8oc4oBXBmFgtF42Ia9wUELwotKrA4NEU6XEx3+Oxx3rwj3qAuCLuTSH3GTor4ZN1
o+gxD1PIe+AEix9xolXU6gsl/S4MbPg2WSK0J2g5Ff/O8TlTEuIl5Ad8k2YShvNVqp24r7DRED8e
s0qPSYV3bP4Rm6Ncyuf1yuSPZcI81JXuuoA2h1fEoZc3JpIZMLRz2wajPE1OzyO6tCmBuJ9ujRUq
7eyXqfgvSt8f4iBrtqDhsJL/hT2fDp1zWG2gIArJELwJFI96vCGjE4TN805/GtAWNGRed1SwGd4X
LSKYB4kCpuLupFqt7BECKPd5W9Gln4dg7Z5/Z+7uC38UyfxS2toz6FudPpVq7TSNL9ehUBtPN26b
fZWPNUUr00ZFJSQ/7Zab9efefQ976y7xUS7Ie2dYYqODHCndWd63MstPFBOJOVC14qaDEvc1Eg/c
WKNOszy3Hjz48pnJ8Gz746aZJArb2yvK3Gv3lZXOo0aTYkiy65NsuI/+GUnpIZuWAw85Ury3FYsB
8abgvAbR+5G+rwnvX4sMCxYcH0UZaLdbcccYLxqbOAWbzMi6vUw8QVKL+qJjYDFkVY8ue3eh0TuN
1SKkPu2gWvYVpJcoTLc5ZV4Qufa4dASnrqmUxEYZZTrIIZPDTGAAkbwciZxU36SMrsjBA/ng70IY
rcsXoGniYtPo0pKAf3Ll6dfltQkMHr59KIFUN4i66fx+iplHsmYJOEcpgyX+W/dEVZJpF2q973t6
RssYJewv9254kS9lmlLBJoM3sCs3ABhaWEpsXL5zc/BG8LalxSPT9hTwn+Y9NYJaEyp057fXsb9l
f/CgnF/vma71/4TVU8YJyWe/b+CMR9IRqWonbRT7KEd4iK6FJt6ZkMqGDMGLDEY8EmdNj5sXtwDN
m75lfXDUsum6N3jsNbarVDnwC1o8sJZmsrROvo0Q+qvozvI6GL4tlEnKGfIl5Ip/5Nl3PUjBGvGk
taCEsBMgS7ZEiCuKYKWca4gs2WyE6Iuw1/PocaAHrvFiAdtTAyVheZ2eM6VPGXEJgxZYYW4j0pn3
M/w4bHxl4B3qXiEFFP81sEOT9BDmk4/zLE/47NOO/ct3NHprnwH9dhJi/k7IU63UqwVfuMMnZUZC
WALxlvme/eaHo2tAE8vS1A4Je7v0TqGokUnl+9IXbpnZgz9E3xEeVqWDwYNKm0AqJ3VjT89jDIgt
F5MV5RV6TFEVclDEHK25QLnlAJpfFC72NTopI/kphjqLeWjJRRkVtKGidwnxPnRnOFdg9km1w022
le3YJh8A75UAIPI6EythBEHXzC8lvFMDs4Z+JEFpq1DYHUsf23+wAuPDrrhPT+AzRXIfkzHnVXC0
jhaY6puG4B1o5TEhz+6g+OBQe+K4g3WwusppQCLN51dDEqOg17gwVwS8//0tmkOCV58oz9KjoAqE
Hr9IrE6PzC1pWYdZi5lfPETAhexfIVnMxmUUbrX3fZaV3OUDJJzxv5vkNneMgYtzhLNSo83ltRgH
r/PWIoTjh+b9zFDpDNxrDZpNQKYPnv9ZLXMBTvGPYniaxWh/ezSbozrk0dE4FRinHVIKZw5trLpN
OcT+g5KuOKH9TXyaFxpQChS9Cw3DVMCGwzCldPojIlptM15f63YjPawqZ8U0cmoPSjI0FdLCi8gB
WBJDIb/uz/nOrx1D7wEQdb0+GA1Id6u0LkJYmZ4T/N83Qf4Gqcxv1nwdiWleZ1V1U7mwswEYqXqk
lmMpgt5bjxDc4AtrGCBz+ELR1EvYyhqCalTCKi95m3anFOkdw9keMMv4tOsdzJOCCN8rFbaL8f//
ThF0yx173Dr1sNCTntDVSwkgGq3NM49PFmSHyO4w8b3LxLqCgRgIMny0vpFVtaaTicot1jgVQhNo
u87QFuKhx7sscGNj4hfPtR7MmhKS8hvFls4CVERpdtITj32PCc8UHtCFGov6/IFK8frhdCh2zXCS
hn/hVXenSEjuSoZWUTMkR0btJpZgyGQ0RBxn/ZRIwydLWE6wi+m6x/8+Z336eJG/POJy/GbZPyrb
IfevsrRMa/NxUinOs+rlek1QI1zwG7DGXr29yavXPnx5xZTf2qhPXKNpyafxtBRpRLFRuUqPaD3X
GrOmhA2uRn0RnJLAuGijlUBMsWNLKV9I9Gh2M5UP2JJ4VlsSW7bytw1EWZWKdpkKMsG2mEoK79xG
ktnxOb7EF5VJKrnNiIQkdNBgubTjlg9odXuiCzWB0OIq/NaxIXkpVlGmq4bSOeE75FAbE913+Mzj
FzS3QX6bi5vTO/k+OrNPf16prkx2vIFjjPjWufMXb23tPVmo8OBl/O2+Fs5e/nIVXpgweSaQZaZt
AbDvyxLsMwZblu+1o4XGk7VTLvTW+BBkdunqYUNV8l2uke0193DUv+oz4c29s8UIZYXEULsozVWx
8m0xEksWcGvszE23Zf7ZRI1CUw1MvTfetj4MS5TLPjNgDx4Btmoy5K+9WwKZFb4xu3j6+Pd5arjv
uS1M/z3mV0sgtP4FyNGIpkYspsSejbBx67XRSBvAQP9QXfGyuL9MR8zUqn2LktsTf1MEmtuY0ACr
tdGlMlx/adiU9OakqqYB013ioX/RnqvOitjXTWP82jN83WAe5241Vqzu3KfkcJpmcS710bNatYQF
EAH+AonuvQsDrUkQSi709BLam6X3omSyowPb2kkC7WQ33r5elRHWO6aW1EE68MLuOP3boDKsiIZE
/VDqNut+Krg6O2LPmdvR3CCb5Q7PI3gYH7yyX9iyIoN1RN7XN9H00xynDj+Co95eFmKzg0Fc+Ap1
IckpvgHeACPzq5jZUlXyh4s4OjHQ5XWNJ6AvVbCcnS+Q3y5bOSOJV7lr57rpoNNohElQUmcSXAVd
BlCLsy/2c7rsTt7AnSYjkkve0m5uCTg6W0jWjMRuquSe0dGbU11bnLyUm0ltrQnZ6lt3iU8t0GOo
3My3PspwcAugTHGWIHUcDW+ztP6olUZC5HDmLcm+TR+MjF1s/9eMf64i8z4zd/kT3WIB+sKOAO3W
Z/8OrJ5ACp6G9RbrJ4jztjykBnPw8k2xvZzJukRCknzRFulG+pzKJj/jDBx1hlvFnh9bqTBTCbCj
1ExZNjj3CWvMDTmV63C9O3d5yk7OMFDz13rDt00vY64P4dXl4HjQi9Fi41DyV2C6/FPqzBvJUxJK
KVCAMFxp8Y09tZGwsvvTnXOemia4EuxA1OBmWKErY8GCPewjCxn+k3yXZOZkmeS/qLPkcKYFtUHx
UraJj4qfQgw1TwCMyfVUHNSw8HwMkAhuk/Uu9vyuyKEDzGOUviGEgA/25jPsdqgtjvXxPTp85r+t
qW1QyIxX1gOzT/5Y6mrEjW3srd3w0zy/1DQONmAdzAof+ktsmrytSz2VD6Gq1OI3LVTGvH2V0iQy
qiTAlCrAdc5FYKbsJ8O0sFxU8IaUlSoarygQdd7EwoYfDcBwE4MohiXSINwL34K2mmTQTbKDtju+
WEHBUHnp8ygs4a4WdZSsvfjkfth3pkMevUu8g1ujhB/tulgpdNVxM6kkq39ftxSf3RYFzXwMeMM7
R8MVWB90GTA/utHD/fdAtUTddxEYpPdSS3aKIMYMHKNrPA9BhV5PNzwTJy4lr2KvCel8jDG6J7R4
AcpKhjaw6MtTD6ZdRFB99S0YZw0Bul25QuZ/nk88sOz4baSCovUb+jqxn1biPCgIHYQZl9A3xmfb
Kj1d+QEvqDQafp6gV4q5juij/yZGrSStJZZrgECMLEFd+OJOpCb3X7Fspde9yr2TWngFbqYfqK5A
H/0hQr8h6amj/RXqi9/M5j2GDecX8m9gvPHXwBMVVMMGJazVkS5NkOLL3wSSjpGuc1U4xlF5ckVF
QhnJwXDVNKPNLl0JzQWwqzWYAwrIXe8js4Jfan4wSdC+/Jw6CKyrd6ionMKooPr725SZW3Dp2uxQ
QD0M3pnOf9XTJgVI//YZVhaRG1dBpFVHWB3/ZGNxGjS/2Ad93AuoVrrcrDoqrAoTMKPWrQRhHdVg
bX27QGvb7cqjSSjm1X3/UrDdvgolEDXiSY7oLnGUUdeuQPeb1CndWW6hGleOsyMynxm7Fhgv585M
Wu4gys5WU5hIOGBNF/uNOJkT51lJ7YmvUdCegnq1l5xgwjPuZCdFWBKvT1bhJVProVfCfLuDpNK/
UFsLdaBWjYJxC6WaXwt2HuoT01Z1FYNLXCp7iQWJuXvUPV6co0HfYgrVtj4baPzNPetcD7YTQ3x6
TS5Vsrug6Z8SdMpTKt/xHFTRygK+NNl2AuCIh9ZvTuaTjMn9RWYVnPPeQZaLF9oHayJ5dJ1GfgBo
bRG2qALy6VoiQ2LUURKm/rhx/wdZ/8wqmyT6siVpB2mvczKzOZ0RBu46cz0m+GOHUXOCenCA1yL1
nufruRVynOodp7H8JQB/CbPdT5U7+KLhrUl+i9fRvzurN/r364WQpvPPAZu5T3H056+tuQpdu/ie
2X3Z5JNT99eortaOJObRaEZC3mRmSZIOZDdyvm0fnZWlA611LAaGZz46Oh4f8nRlg6G1SjkKaNAY
nVaD6dYyZajwiWQ28o9Mapiuo4S4q7bIMc9xkuFTe6ppmJifojbE2KmBWW9i/oS35L3rbN37qgDB
7Ul62tsH41gP85eCG1MimqJOIcOzTsldtHPnrcN34QSDcR2oP3Q8nZgYIwJkBjOTJj0WavcT26hP
TPNp8cQmrP/OOeC6u8MkxkeGjl3mDgRxKy4N5URPzFExHuImfU9cIymFTIWLSHVqTPZIERwNS09+
BPbP+lJiOdNgbyiSduHBNftbWRCG7cdR+1NhqfZPIRq8B+snow2AW81AevtQATZi0P00NeHQ0Xsw
5Z5DFjBd/K49heQZ3wdpxOj9+OmuQmT6i9jC6YyDdgaYgeeari1utpMFDNHrD63NnqwsEyJm7jVJ
woN7BsMeqU15lVJ1o5JeB69nGJNmW5aA7ssy5SGQgidwqTT2HMcqlQsbLKTjfSzlZfa3PoHix8qK
I6FgxRSKObSyyyAACyYZKthC1UpCWVEIx+imUVxCFea3Z8uNW/U7cX1JqfJtTeF9UmPWcrCV2Dlf
e2Ma4aVKwJokoheiUi61DHg90s/PoXlz4p8gHhn4aZ4vVmFCzuugt7jDWqxb4IxQBLZk/CDj5Wg2
NQQWBUcZXAQofM4v9Cgnq6GmGy6L5G7HtRIzAn2jTh1BWjxqkuyYNMS7K1psqJoZcO/yXvsGwLCr
QTkffHJ/pFzcQq0OYet3FjIZuu0DCLgBsTvVFaArFomfQ3PBXJff08f2p7HDijsZ3EQAFR8RPq5H
GQrn4G4iWPVpNL9K+O7IlqrmuNbg3tXo3U1INCJgHAa6lFMnFdT0oIwDwy36s947NidX7rfF7BGF
Qzvy3Y12J3q7adr5WQpsTCRRSvrcNP6g6XdVOUwgOZ32cGXgaz3y+fCVPLqLhhpp6MVP7lXi3i1S
KtQOMWapEMKyt2zZXmmr0JxJBt88fgSIVq6MT0+FYgbxAHdTDkxGwkNbhEd9MliKhbPw1A3Legra
BquUXzr2qKYl/AFVfaqa6YTAnWcV5JhusSNEaVWY4Q+UPS+9x6SLvCiHnGdjlVQ2VJqkn1ikSOUF
poQUcblMe1O5t3FCQwMr7xXKx5JPGdqaP1dGCuWpe0GZ7y0iVPzBEXz5RJVc4IrrJZTz4NdNQftq
U108s1pvr0Mqi0y8OJvA7gSqqijjVqjEA+2nxLuNsLJTHQ+rfzBjLyEqjQs83QxrTY+luW4CGb+P
z0y2azGGFAIhyhFgpUQ843QF8j141wUMYHPuXLmWe2MMTheC2XyqTAyDtdpdLk4UZ1cpwLb71b0z
X6ACALT3c5tdK5lOWXozsTix0uQjKNaNxz5jik3rFElst/kf1PJOW0EjxvQkMKVOGA9Ww7fPHxbd
0EMITeb5NEhJ0gXvbmDgHLO8/aBILqxRRm6YVwKo9AwS3KMkV+rG/kfubtGJP2EpOnyk74SiqbEI
Byyuxa1zCqKEsdEGkabjOV60JvfNFuqmhui7uIoNXZeqSsBCeHCNj7ap4Sd0F/r1cnUX5Wcu/yKK
WnI9I/SHUMBlMzylQvV8ybiPMJIOs/R8Rb2t4qzzSwsBzy9N1p7MmFmkB9dclqlewI5IqcZo9mCS
RVqqSNbfsNWgHepNv1NyR28sdPbyPKs8SEkVfzNEDfvyePHN8x6Fj8C5M36jK6rhiySoRmQ/mqLa
ehPdWUbZe99tNMHwOA1JGoaSpjmZVGQuclfW0itpWSkNTyGPWkMFKNj8/RPj0VYNgTUv3qdoJ7Po
jYuH6rs9dgCDL9a3/C3FBBthqcHntA9pPplrMOSeaETiEtfJOSh20qG345PYgAZrrNkLjtyOXwPD
Jt6D/Gb8Cz2LnO84EM04G7Mg3KXfEjalY3rWP13YMrb2bkUVG2P0f1IW9EfU+JyYuLaOPkMX0o2G
LsGzeJomycY3imgZOVCPIVoXc/+WWYz0P8MYEybLuaXzVhlMH4p5esY1vT2Tm/WlQ1Rc8AHuwrr5
3mylqN0ymNMaxRF852v41riqTXRIoGBcUSHTvonOQDJ65kTC/ue8s1V+kDKEnYR3KXZGASEp6WLj
mK4HX5cXsf8CZnXbQ3u5dLfpvBjmugTo+nzfXtDr/rMrgJ5bPjGiLTFyn0peCf9/pGUyoP4+l0tE
XST8Ke3uExf7OisYEGseVTkSz69gC+djoVwqdKA6Ipz69WKmoqCj0xs2KXh18EvRLf5Qz/VKY5MZ
UsiuSAtZ0qh98IMZ2M3ls6MtvQToS14Txq46Wut4P2pPGnb8wELfPYNfgYJacNg8l/CVFgE17ZZ5
uMby7c+RVBtQeHrPxviPnBLHgCp6vXBFRI2LBlSmWM3Pmp8qn0MZYf0ION82EQ4EyA2bGpMKUQ8c
pTQBRVaEZ0cGBN2eGhk0b5Gl0iDp8Kqj71dMoSTWYghgnaAyCg7+6mXuC5ROKXa58q1ox6H8Ux1r
qc/WsHztyeEKxm3Ubp4sCmn8FSypELHHYeAh5YhRIrXktNl+02H7JQbb+ksmCli8tyLcbBtLFRnw
ujMezces4Tegn4B0P+oemxFlOOShrDirAV+PxUr5189NyxhMElSrFhdj41NvKp0puB96ue8AnFy0
G92YdjB28qOiTVbQkZxlMxiwP5UoxhGLMpeb+pZtNXPc1RobKs0H4PRV4ZuD7k5eqPX4/BY1NppR
oU5gmzXR90xrJtZuLLClU5q64e0g4ystli86kmwlCiTRygAAriWmToFa92DLpVPnc8XIfX9dpqLb
BSxuJayZgSt4YanVOsFPu54SqE4jjqDnPbCcSqCGgOGEQeVnTPt52h9+IcNsES8jUo/LTvhloqoV
JVconoagG4nymrAel4+v1I8ppqlBv8spamE+RAOxoXIW/6oOBZcjlPbZpt2JB/AUTAB3GLHZ0n1T
Hy9aApiz4yeGgZVdjWHb2r6CHBdMbNKhR8Ri6APoO2gfUaHsym59eGxrt3rWl9SEQU2LmfOJsQWi
3FdK+3Hy1k4nSbiyXJl36dwt/bxy5iQfL6Ax/QkzD3cDVkvsIzy/coCsKhK5cgMdjtxXmSyqcmPC
4pFVwZIJoGsBsOAn4SbcX088yNLurvjJrZqIKoD9Y+lKdilINBB4mcU833LXMgOrPNvh3KmJehmm
blcCmDwMLvQy3jQqBE9nDvO26H9PcnL+ypC4nJqU0YQZaSuY7+oXKJJJKBgGXfDC95ELNMKcxSCO
6warMlvIVgOg6ma4KfW+eultmc+6s1aY4H81O9ML1udYZW6iDA6OXliSKgCA5SrfpjSHIFKvZRn5
csAdWEiRY3n1vg/AlFuV+GS0Govnh4/vVmKBYHulUzbjwzvLwN8tfy1XZG3hUvmxu9D3L6Jf2jiM
GxZld9IXhyiPmnukUF+RC2TpWMn8m6gRRx4qRYSDozDR/18tl0N0FnyLE2BwEACKqY3tniZt1oBy
nFTZrds3fYYgBn3yCsDJJBwPJOKDTCH1nIzIAif6GBfbWvy1UbJC48MX5Gtg05vm8UMLr4tio7xf
FVML4EhUnl69K8aeU8BbkVBRHRor46bqBj9SiK4Fs9MYNuxrhz1C0OJQ3ViXt4Ztbr0F5Rarib28
C4cpgoPt1R/CfZvJtX/1txg5dfrT/NeqfsUTvT9U003RKcs8hFfTTYCYLCNJNsCoCiMqPTr/HvLs
TTUGVkIqupHx+RkN4YI+JvWt/q8CDDZgoamWgUrJX/tQktdYHG96uBhFqUsWAlLEnWDXG5qgLCZS
Rca/dS8u+OAGgOdutUBKZtNpoj4ZDbFY2VTsB7DZVXm1tyMlrvdIglvhX9WsWmXypmaBxmPkSgOy
1MkWIFXF3t9CvtahM24eChspxRKsw2WI9uI30XnJg0IG/99soLbK7K5/GY6KSzyNxo4oqwjvGrkl
BHqXKChooPSdz37T7fJHJjqsjplb18QqMswrSiuHSFb2y4JGpL9qT/p65OgXhcXsORgm37oO/0Th
+ppUETl4ogNpVyECpRrAapmCF/FLnfgecwCgorSTbhIgh4tFzQ8ZlebX0G279AgfXStiCmF95nN1
ZFZ4hO8rsppOjAJ0r61mIwPImmBzr5uh5ss6QpjKCu6j4a+dGRv8GUpU9spzBjGlwwC5IIlvWXkw
5c15H86K5n8C4Q4zEtfVkrS6TN80UIGFGOfT/CBCaCiVnkPLk9l4L0cpYrv4/9hBxBRPRq8xoK5K
QWQNy2AZwsat1gLdpqgnkneJW6DW9ntF69uLO93LkZNJc4YCdvvUNP9/bUINX2cBEyXuGlthvUMZ
ysRfMSzUHIUUiGntq73O0wE9csR411IjFtTpD76hQj0/sXEclSlx9wm8FISOkXCkWdGaJx7kTG5g
veUZLWcZy9gGGnToBj8Yi13OCSP7IEduuLtwb0t1z2V28HCx73BkiDMrhsBOrPtwDd+mLlbY1MMM
wJ9zBRnPDLlxfSotuGBoNg8l/gTitK9jouS7MC5adi0Ek5w3UWkdRgz3+X8FfM08+RfBSSjLt7fO
S+5o2tBf/wHnNDx6mSARlGfYtgmJE0bSc6qwyQnSqrkTk2sNB4lhIR0T+u5psNRJ5hDu5G4StSoS
lZuiPPVIIKz75xoRbSgPwD48c5Xp/6u0dexVWue2qEc3RwL8fHMaoygm5yzdOwvVTCbnrQKHo0Fo
E/iV8JeRCWSPlOM5EQH8Bhf5YDl235dXBhxCQf+BiPeH4vKA2UaD7d4WRsCkC4Yft8+zN35oGQaO
7h9ePMtDB9wKpFbs67SfYt9JqAMxnBLydJgafj/rGTd3qxnEmEueB20QbY2Jr2pybvRS6g9vp6JO
0aZP+nVJd1pPTl1GSAtmYmRvpbz3Uxu44fDL7mb22vHz0C9Ow+dki6GnXr5TiCYcKqMkmCSCRua2
BHWpkV50j7I+1qHOV1J43rB1eX31p6EUb4F3zY9vTMt96ABToYGfGlQliWSkYkpo0DIblSBOBFUw
YAhzsHKx4u3c8Gc/ZJtJE7pmsW7t/jlaNAAHXP+iAM9QN4CYvEUiEg1j3gSZ2EwqRUszYfk6RFC2
4n203JhkAtH93CndnZpxmKy1jnAknr6ALf1kEBKLXJ+iBvKRz+VJfqXJf6kOi7GyxdrqSph0Qahm
fMJayuSVXcJ8Z3eMDMo9SSQhszSxH2Nx6VlH/vNZ6gqV/IvtY6l/EXkuFGTdeOSG18P0hLFRW5qW
1BrMMLo5Gk8IPdu6yVvxGMevC5OaMyLL+AmnwJnYj/qgW8Od6xGEs7K4d2+J5VeGBnqRyV/FNLMD
uC/g/ebwKBWN9yqDKf1CzKx1s/jQWn1eBCV2kY6t+xPvnDQill4hmX+SaqJmG1flhYtxo8rGmWjn
qw5lAsla5f3JFa0ya22feIdSSKFR8MDrC9CtN5W+MLhQdfjZ/3gLrxo3fDLUUTJ0uRrGnSaKPo22
0Fa7ROxv2NyBMvQa8ILytDtBqdWz/2wlHBJ9RbkL3AQ4GJ8bUWu+Ykj77grtIxSMm78xgcvbEQH4
TdFRbmRL9oUfXrNpb9YHZwz28pc1JKALQYdsRmttl9Hm4AIvN/YSBhdO6rjipPbRPp4vSIw9lIRZ
R17rTh1zYz/QoCvO0EJkD/JfcXPamDVDu+oh1hVscC/djscojjOwPRKFAimkNPDdmCLhZL/pCyA8
fnIbq4S6DmkpBCQuXgRmKF1jvP2FEXxjUOKZhEr+luw5RRbRVtXNIA4OpjzUJsP8rK2I3oJljz1B
yOlJcHlp0qlNmKjQBuuj3Ag3uIh7NDRhmmp1Vcib8MmV9Sf8blyGQlM+uGp0izAbxOdcPTOurc6a
1wbZV7wBPtHsMBuGDXlYl6bKBH7Yh2j30B43VvZJhLBnC99I6yr6btb7Xq9ZkJpKy9JWnGKIUhs4
w8vJV7hiISp954tAJf81oVoQKcNBw/vn/uc31lfypqglBdp1bf0vmvRSmbEauP+WZHlo93uKknfS
ekRS+VAl2MfKnChNxJ8SPsClLRa75HR4XizRcC8vI5baOf/CaJdj3OxxnAgGX9VW8kXZcxBkdn6Y
b89mYt8Q+wFzx3/z9bKd5mSHXc9kmJpJQpnFRhFWfUvHYCrb/lHXo8FHN1LyzmQouYC761Uq9M9R
V0gt3HbgrGWxlTnDctHUyHbLhj/zFtRjragAbGJf9NGJHZ1pBFuej3RXWSEqm2N/GvrG/dmdPmtx
Dq/v2zaOu+U0k27m+LkKCWuT4hsx/lZK4oRKdFPav2ZWgDzabYWF7tkItmiYXG94hvl2SPHpqPZH
yWgka+24I4H2/hhfTdyK0KpQx3VLIsgZrFCCOYJai9EdXonDN+EALjkbLAf/190eaGuapIpg950O
GbqQ9x8MsKihTstKBB42uRtZOzZoD+wVdVVgITmiCSYLJVuETed2BI9lpmFJYLLY8QMdpAXEBBLp
ildfG/12lkRo+SaJMfPOMXbOp2IBZHR8zpJN84llXXtVb2X3VDgoNYCw9SMgtRmilWCRUcHf8inj
3Uf0gdnUH7P6GBBKILBM5A1cwy2hUoydSjPSdaYtUFll9sxBiE31eHgthJ5YQoIngtwxa4pBnGYH
alUtKSplA4AY1wJrJjwvBNwEL45fIqtU+G0ApkX5qSccskwWjG/fqIgMba0Ff0ZNSYCsx5SkKejh
F/8V/zgq4b34ASlgbKIdlxlPTOzcCGiLvF67qC7YjiEHYEFGsGP2mrh4aK7uCkVBfSNAe7e+7cjV
AaMrzgHXsvJwsIB3FmM0aY0QLwhEHP8TcbGeJl7YE//OHqjY4a2QSSxlJnizqqARjypy81Czl1l1
MgYGvMwjG7h3TJ/ljDpa0z81OJYL6uD0W4XD9SnQIEO4aIUvMwy3DGJJGfpMgpxksH2f+Jkkwsxu
/Ggbpiz4NBXMe0YhSiu1y+qtUM1VgLs45ZawlnLEMuj47h0HuZM0ww3BOPGaIgaNB8xGWTIdS/r0
glk3tQhVYtGeokEr76cAgvpMva07iEP6J4QH3juCe2h6FBzlXO+dy3L9T53XxDFIhnS2iSRMtQ6Q
WW964ji1f+ILNEnhEmD1clzk3A78cZ2UpUo1FlHnhd1BGvm4LttKLMH324jwR6ibUidCnANS+EWX
38fDuFUxLpRpUz2ih7zWMahobwDQedAj8muN7jojrhCHGdVM1ezL5dH7fI2BWOsw0zhTz96AOsWg
FASyJIawkJvWf9toDMEbZN1Yhokr7H0SM1paMf7XSOkwowr+seH6TYUhDSzbMkNayypt3fjrD654
jXiWvZrN+xB7v0KSVhiaxlVgWgHFIAKDcOmaW1dQ1NUYbSjty1GwPYWsO8DVuos08GGFlVWSjHgq
6iBMn6tIVeoBnxPiPuykMgjBQRmkJHLubxojeDlmGLFTM3TfcbVDZ2pW9CruzW8GHC62hF9uwepj
2C6L+N3zS+jM6Eg7mMyNJfKpNmUEI83RGnGz5Nihlr9c6QdGeOlU8/Xsi5Hy1BPg5uNH5Xy20DVx
nM2tvcTJ/C2N4X3WI7NCjWGRVSuCuhiB0xPvMzqJ1z8cZZxPPqIzWIFMVJuehazkLlsgc4+u7D3e
aYLmcGeM/OtJRqW8spHQJxFiZE4n36boB+6Qrn6wuYiib7JIfVzKY+r+x0tcwupjTUTiBLqCt1rx
CeX4AGkYT/MEWGwTOHjFoazK0gFIQC48X74+OHeaAxWxZEzK1kwJpIjPd9SXdbZLg2t1TfDeQAWs
XbaLjGPoAGZQnyo+HiPcHCDq4Q8mQyJBpzRyyNvEBqXy+EnQKed3kjER7IBDBeg2WsRZ0Mfgg1mC
0IzjrWlty8DWWavwIAmOtTbQdco5dv/ivGzmi3pgSCq8ouI0VYewCmw0h8bKBIswTehnIcXY+0dV
00GdDCg3e7H7SLM0gBh5DyrwL6FH/9GHd9zrGy7/B5eJA7ZBW+c3mIf4H98Bq6GtSiTEgo3DMOZ1
tAHY4MpH9Rdi1GFBg+2f0DorHAxtkG2OPk9DN/9Jai3Jz9qceVRvfD4fstHtf1X+K8quEnOlzEOc
pS7W6ff4MdOp4QMjTFyb2E7etE8upbba0CcZmSbfcAFbb0dEphkog+GmlppyBm2dgjvMDSb1c22C
xQ1v4fEEvvFZTWsHfAxRpSY6+3mBbNU9qsKwBZELQfHvyvf6Qgf7IWc9R3x+doVGo0yathLtMmzO
/YNMpQsfPUYjy6jDrWjo/XX5BilpttwCQdWX5+0QqJZbbAnDv4i+n+/VFyGJvo+418RwOwwLhHDO
O/VlfOk1VjQLA6ar6ClX1xh/IsVi/Rwaj945gQH0S66eOnNSJ9Nit4b+A1JJ9PYRt7Ieen13+031
qYQscKtzD8uftdvNfkygh4cGpbgZ6GoYAh7IzJ9jdN9awre/z9XvCIqjTspwSL6rBPjgB15jFRhh
emVr1W9PT2Uf0gCpE34QKqBwLhRxHEbR2reVqOrIVSsKLryGVrN5RM0KsY5O1tr2b6T1p7Q1tUfa
GQ0hA9tcL6II6Y3Z6xohWQBAr9TfdfupWJh2QuX1vh/2sHyxRSQLwK1xKIcBy7O35qik2ivk0/Bn
eQl9D8qjH8j+TpDIbg5qWgQ2zKAMQO7zI9omnPd6Gc8UKG7yVGH+nDHccwATCLM4RghpKNWJZLLE
gpx7Y7H29eXB4UhY0akD32cFLrsKjbCHA07DAKQ0e15/xXIInHvAMrdn5UqLnnmvwnVULZC726E5
eFiCnix0nEp00AHNWbx20+tWAw8qj8wQdgVTR9MqqTaO1a0kvriXxFVf0Oqjfo95JAuQKLPHDfd5
BZXBhk35q5XEYKiTtFR9GdNCoDtqcgdoUzCwQUiSG68S+VMrMFDoRr1nbUVOaTF4XZwnXig2dJUn
JKczIjWDqfsTCDu8n0hH5hMadZV6SoGah3ww0VDlCGR+KfdYddY58WQlcS2m1fFjl6OlYBWenu42
51sIh19yeYHJ13rMlZNAd3yx7INY0OD0AjZ+7HyebKd8YNTOHfVQxaodK9oFGW8o632XHewD+FUQ
59zO3f006zFEGIE/1Ixer55l4BnwcoQHQu6TXMJpd0bIpyx/R9niJ6XKOxHqO2krgSk7LAS94dZ1
GS6PjWywe53JP73Jtovs7MttE7sJWqBBZA5pQ7gF4hJxWlqiiKNWALA2CAgTaqMWyUeh8ZZIoncV
/ErZSh2DWU4cVrcdmedNtOE2AKrGNyg/Gw9c9MTG3hypp2STu4fmyQEyeCq1aZ+Jhy5VCybcV+tA
oFhoA91nviV/3RW0cbNWY9+W+uQT8idS6MWmtoOvoKmE1r88FbLcoaYPyApWFTQAEt5ggmIM7u+B
u/ckkCuIvEu19Vm39fVo+HToazjq5FML0tHDgcZhpvf4Sf48Qq6ONLd038cCt4cnLoV1SPp/6ajP
E9l7yRsyXFeo+Y52TdIizic2pSFIHBp1/lUDe2ars0AQdnuDIa0UWW5Rq6qA0fc5E2zzsVybn0Js
lho7rg+oENWV0FncjPiHyaJXI9kvNpkmAcY8JDTi+5NQ5OAvjGYAdcECMyXG7AD953NmdsslHpmf
pFQ9AXMaa5zQi1WuG7b2U9og+zHHQ8ynV01bzIx7Bwz652jKR7gl7FOdcBKyToSvFu5l9+ZqL387
xppp8rAt7Gh9fErBju7Qt+GxorqnfPv3cqqSz5vgjLI/zRguYrSW3W2YvZTXXg88MYCL9VeEoISs
SCRBmMdl13/qCRlkTx8ewg+ynslNSfRJcDA34oUw8qVr5QnzZ+HqopCv1i7OeMLQmIMU+Yhj6kMl
DEEaAt9QI7zqYc8iFdD5NZ4OetDwnRwu4yoh+q/aHV0REOGrkk4hTDChKPGIRv2MovR3XIYgyEle
wEXt+LOPp6DEBm9Q6pwvKYYJe4/xUkqGRYimH3WiGlmtLn9OJmjynWii0ZyZw6RcqRwjQegMCJ+2
LI5/wRMBY9Oym4KPjyD6F3p8DZa35VaFk5m1O7kWtkgXYFzXEyP00JDM/yMkUKUhpzyv+ZLVHCaV
eq4xluoKhA4TlOzjSNVU5wetzrK6PMbHKERxxAhi36Se3jHDrzf30GMoIrapaHnkhMgy9QX5pcKp
R4UKq1K9txRNSCMAJVLpe7aqkHODKNyQLlC7RbhQ4uGAdK59dOqMZ9UA/wnwKIvnN+cdFbSQjIGK
EwcypGT1SCcXbuMQU1OW2p5s3SCBqZZ024p96neZu/PszjA8rZeMlrijEYIjuP9Mzaywo6xZCaqh
MUB2OuVv7KOzlpswU3h1KXhVOhKnY17MtSTFPxFu2WVFhr9atAKBD6iA/1632ZhjsQjkzQhwVC+l
H+rOd3HpmJrbsuIRuVsEzpCkp3PcsBrpalwm6izGl30kuAmPN4+a8L7ZBKkiK243F2sDLXIjiD0h
yIIL0KpFFIevhlZaj27ZOok28L45r9ZyHlwc48ZJDNfJOjJdXMv+nPOdv8D2RbSi8V6LD9Ylg3SP
5jHG+hDO+xxgqbOTR2DjIQ5/a6SZlnY66up4d18K+AUSXtYFfdpxlhhzqtID+mG+aWhtfwB/3/g9
UNPD2smDpECtFpdWc2pGEo3bOXvFGQMatqi6LuKQ9epvod4zfZCli3JjVwHKSGtuH3nAvD8CZig0
F2lzgtS1qVYndxvHEVHg5lgJyvHGlRA12wnQKAYN7gFoKta+Nxx8lLgCBq6NqyjVs4/zuTS1RRjq
gIh3RrcllUSZF98sw1wMalAOxPOY9FnopsBRWEpEhrx7sGe1U+tnwnksdX+RKbiy7zpJExedVmPq
tmSwy8G9HyAJCzDngrE4kLRSLb+RuSzOOMsNIpjTDIAf21pwqTQUKImCWcao1aH7NWa8npiZvVnU
7LDq7Gaz35b/H0R8b84mjgoH1DcEb5DfFsdvJYc+1ODZ9tk37CAHGxuuswmHpDSM3dqUUkC0iZOQ
EIMFxnbDJPfuGUgi0dsEshmdlsLZbNsC/zYHVFX8Zw6BqElqI91VQe7ojn8LgbzoVA1DhHjBkJEb
4PKkacPe7nOW6bF8Y9CmhHxIdHwgbkTyKXeBm1vYZlBujNWiIgxN2t2t9wzUT4iL3cbptr/UeX2A
vBcsjqKhMBpgwBeSUor0eRFsWegbEM0Am6Iz/OQRfQOvO6Wzd5SO7812Kd0poxgu1Q6iudmxMKHU
yeyacKLKNWbA7cn9lq2Qg4IxAogQ+C4BRjaZUcJRxw4RaYlzItevzpuGf3JzKt/EZWjFKeDsnFsx
R0a3FGrgMz6wudADXyS5tVEsp56RZRoUeVRXXMwauv/gnncn1DlVADBS4cJZ+evNN/AGOLxxANNd
EnTNxI/4gRBDRwcBijCo39Y6SIOb+OocqjfcBse5/+RWMLmqwJrYAwgdFIUasxnPM1QVkDQS9n9r
g8R3ogSlfGS1FusM8Do3nm7W8Afanemg8LnrWr+e5K00nT8XiA2BnOvEu45RBHgfIWOEb/pJI8G7
QXympzO98/dEXi/9VmtS608YfVBxZ+1Di6s+OwQtVt2P3a9N4Ow3dbFmhxrdHEfa+9MHzb+LKtzm
s/N4Kzjch+/fd32Nz1yOiQOUdtXboj2WuOw41Co+VEHj9KFW3RIuGWqIlJwVOF0lPiKtbXJ4yl/G
jrSk7PusZ19PsPPTJWOXo4eto7RUJwK3tCJEkH5L9WV9eZnCNW4dmh0xktueoSjEVyYiv4fNy5Ce
orqueCQYJiiMDDPk8QhyIIOHHPvHU7hpAhJFNjbAZDmmj3pLWxSH+I2PFzVFhMBArILI8BmiRhw0
hmXjGJLdz3QbKlw+g9GisZtZUQq3WbhiEkcljq6AsgtjjwYIBRgjMldA8BixHbTwGCljG+wutgEr
4cNEx29iaK6M2Qgk0/Yy5jivAsnT6z1bjadS8C0fUuZYJ4JoPrbvtZk67aH/T3lepNRJx8dvbkqh
z2NM/cEp7bO/F6s8qdF+kbZZwIrAyzX13Rhq6YsISC9+SnYcYlGQrvUUtFlWLP0qFYp7cEoqTF8C
RTc66d1ha29eWtEfegVm0qVkfYAJNY3Z3UlFohXCJCt+OAyNTsDIFZRs7kQ3fAusjtWonMR1AG5t
9n34vWODWYWGmE0Xo3DCMZ67IwyotATNIj/gAyacO9OvAK2RX3nSKyiylIkQ+WbD6C7VGpeC+7MV
Zq1LpG0/WwvQqarO3VyFrZ0cNOuvU8IVBTlRipudBHxjeN9jwHc6VqYb8BUBNcdETHfdFAuX+q2f
XGiypE6F6HhElkO3GrPqaNT6P0oTIaGPv7xnXKHaz+VbMVACwjLbRKqfL5V6nSGTwu0f9mSxkhSq
UkG+SdvERRTQ7gGjhoY7xmS96Hs02LxzfgdHp5JfCf5whrW0W0jQ0ZZmn7dtzzwzs5D5nqT4sEdn
ZgXIKT82Ao3NlyO6mpugR61lQB/BukspXIK0wQ5UbaURMlUuasKo2TO5b6SYP1JdNkda/RhPww2f
rPccylk66/DxDmEChsrZfOBU5JyzIkKEyVxgX3wMvoJAiBoBqS2+uRk/afDOy6dLa+1omCsRWUba
y5MxK9zfECSBSVZa/WgmVG+cbvkwP/8dfoAdzEFjTBCxD9i76F+0DPjc2AiCKmr6GHffbldDXjlR
hi5oPS9fy7eQQzotbT7+m3SE3FUNf8DBPT13eF8TuS7ARZzf8cjsH1QWag4UHie4fJ3qVG/kR/TS
4lQmtgFkg9nrwXimjtAWgabp9a1W5RgAgZDb+d1HIEXE/SUaFq1JliUr2mORX5wjGnD9SsTdvD9m
83qlneyO2goNteRAbQTuctQOUpaToteAoViExYYIcGHUAaQwjp9FcI3jYB7h/ooUM7c2XlBepNgg
U/yK4anI3PExoqzf2HYyQhPlCsHkALyXM9+G9dyL0Zdpb5ie1hCmDeZo1u/nA6LRmIjJUl7kG83q
YYcGPYnnY9txRjXWEJ21gF7uz7CIHiJB2jK1UVfjG3XPjEoXbGtnUlf/h/lJ0YuSvUV6/t8eNkJS
Ar6+sjGxxdBUzU3/UEZKrsHF8/TmhYE/pkMMZxoVFjTcLrhIUNDX9qZWgw/r0eZNx2RAzJP70uBV
Ib8VxQGddOYln3A7VE50mSy8DQetLQu1iZBTIZngwCiG20QM/1yt1ZWoqjRqOI2hbAEe2iklSCQA
rlBr7O8JaWyfoP6BAHRhuQz9N2HijU3kMvrqxKzLpeFNMbTbJg1StowpSXkVWIiG5VAaQqIXdkbe
9AUr7o3Ez2UPwXOhZygWia2xxth5KQNDjTeoPGOufP98C54cDww34p7w720rkyyDc2iiaCB6cipz
c8HPxjORJ5zeJbEhOynHx/7iKun8x8jTBM3sWx+P5cD6kKLHKHLZFlX3J8/d7xCkAEIGHgIK/Sz1
ZYKV7iS8ukHITqO0r7g5ucsyI10bE3HIKd9K5j+GxK1Ii2dwDwyESLDTMhVsjw7Kbx1epJn1hpbk
HHbiv8xE0lEakWGK7Yjr+6TH9oEwMLCD8Pke1zaAYw2iMZOafpkjDH9XnEvqYAIju7JHr/dWX5k8
9eHIkLxyu+cUR3O9t3Zad6ZC7xwquq029Cd7DSSHCWkqlr+0BzDudcG0KkZLX0mf2QEONh7dntD/
n8Z32xw/L4065e2njSe85HQ1vz/kpGYr6EKKbmeD2Qf4WgQASGK22ZlaeN32GvAKOG28cfbsMDjQ
cHKTaj5hdna0AmiTcnx4qLtNwASQhN2zqJ/g3WgXQoOWM/+pKMjCAh/nyG+x4g3SA9C5tXc47zqD
ybIFzFuY6kAedwkCJyEd7/y1yUK891AmgIEYPx5S7aiYpETV0e70iQgPzEslpZa5QegJMBF2+TZB
0kn5cG6P8pnd+hSAvlW6dYnaXNjgXI/5lHqnGyT+a5cuXO/80dZDL7lCmyfBD1OBZmTTLpr+7k21
+OwyH2jiTv9zMyNLxgDx/lX6MQj5oUdchuRiHpntizdW8ef6OtdDEFCnFyFFyEkPHm+7JwFTIof5
wBVcjo1xixwk9eSmmdyHOaPUQgtqMLf9m36KZmjlYl/HTRX0FINCRUCSiS4T5OVD7Ptt/PNueUKr
XOmPltlPv0fxNwfof6Cg8wSovJDI7tcBbt7oViGqh2zMgNaoMMDRh+TbexNLXPR4z15zTS+lr//r
Xa+abhiQVaNKySytKEi8G+Z8zMgbAjTFBC9hb0+Nrg+FQMXthnVgvS739J8jlHd5tSoyKpaX9nrU
fwidsV2yUx5T/As9AM7OuP+OfFXOKHAYmn/IR1JQNhvJhdhXIemoEAZFgNu3syqu/W1mh9ZIRgYy
zfTgW+xmbpGms4DA2ja0fwBmSy++riqJpkvjPFx1BkR0pQVGABRYOcZ4AiAOfImV7Jh6Q+wz13AN
bU2h0ThSJDAVx8lK3SJRW8MfSq6oV4AnCWd1nJYPZ7ideG4L77Vabv9wIU2Dj+1/MJ9QeJnqzmv5
s85jGpbolFgurwBCQFo6a8xO6bUfSJky8ZCXE5ZnffNgTZI+Qq4O9+HaIXBpd+pdKMTb2vUZnNBm
pglkBgXuuT8K+pBvpv9l3AXqwkrV2j6pJzqAhSFfBo+LSaHzgP6wM4HhmSeRYuiF8VFaRTgLPRuJ
vWpKRy/fAjwYgBa8mYreb6rrnMm1/bJTKtfmlSKz5RIMSQZ1Kqi8jbRZT4OvCP2CLXcpbOwVWmGl
0FYB0dHF+R0Jwam6K6R2LL6JyV+BQkbfg6FmuyFfQkz+lPbLjdGNRjV7GNYAQe0MYCA/fh/HnWNY
CpTV6c1o2d+AFyvzsk3KtkJl0WIv9O+KPjS1hXT1xk53nMN7jJ0YBdlnfNkv5fZ4ZkfRG4K04nIj
FMYGw6XBFjbl+jnq2Lj+BRzWEnQHqPIVjaVuLG2AX5sf6VC/obnM7x099sbalvgXw3mERVZV9vgE
ete4icoYASpFeIsdzl912rI8frxj0poUaP/eAs8zBXvBanhhvdJ2Fyx+TD/m8F6AK/SxSDnjhuus
G36XrYJ5dDvHK6kCiR1J87pSQ9TpV6R2B2pRgCTVjt6ZJhQXlBI3WJEM0egF9ERTDIQhOFR+9DJm
aVRX+DGqfyyxYR503jIRzzf0C2i+OE8pSPk4RmUB8VOjUcnGSY6kcKLfVjnLWAtrBZOBPWP1c/Z1
+954FmYYfVyPduHXXESMONpHf3xFys/SGji7i/RdvQPGPOrnMILJAPIk+sTcUhwwrw+IWIJmLWMX
MYm5jpYgCx+aRhY1u+d4bSAjAkBbLg5u4JCtbxI/vzhTUBYKk3W2GIbikXipU8KxWOJYUuw3FQ/x
T3NVMsid7gRburXT74Onhh1UgpCedclgrP9ZAjM9eSXpMo+EurUxnaskCaSdGVd7AoTBSMwlYVph
Af0buX91wMwENyc+k6TIJTvlAR3YcO+/JuOox3P1L05Ah3Hq6OEhq73AG26yWSDhLxTBQ0oyjpQq
oLCA7pAuEihyIWYFtDvwqzg1Xh7RTr1lsROHRYM96CGg6Ysa9DqSVdjrTDSj7KC1sJiPnAFvabyR
35SyvfFy26atEN+PklpvTfNmDJy/lZri9LFd6PuumiDkeaGCf7KC7iLDbulsKf7VlkB0PQdOvTmT
/VDZiDmWTGjL1w727JjUVGAak/jOxczau90OjUet2wLbF09z7xDMZRB4/cJlxQIkPIHl4oPpsBEL
zTvlcIjoheXsdL/ERUOLtuCNTU6bi1QhPnN78/++9EoCUFplE3fjthlmWWMyGaghqNIczwnPtyLV
0fgl7X3dnc2AV4AkusQj9J5wh2iKal8a/EjSbnbwLBmsMdU00vaCR79BCNMtglFbHwXeFi9heQI2
xzcDsfZZzsAGjszUeyqfo/n0NMFm/2ejTmQy9JCmCAkx1lFM+Z3eKDcaUsAVCrbRtwk+bAj3veZ9
lJvCTV6cxpnIZiq2i/oYYPwtY4FJ5DG+qj9XMfi5ofVEPrlAv/RqhOlf7XJ0y11nuebYiXN8CiYH
LGYz6bktSUq78tax3JPtE+gff+iraP15+RKUL9Bv9ngNA/buWrVExrj7G5lcTG7XiyZu/JDZuE08
WTkgAOE+jzg7WhgTiRBBqja+ksFtHZtB+NboRzHGwpIk1zSRwAbqncwmZHEkA4tpXc7wiZ5ejF+R
J9/177eD5/W4dxvBv4xpnE92CEGeGZ2HaLPnJ8PuuvWXqsIFlArNPba145RpPHInQG9bZozudBox
J1QhNRX04kvboXFHlLk3taaUlf05IgV3QKsnse/dBmXBlTeZ8IXL708+M0C+sxUtNqWl6BTLKx/R
AcCz4iQurjhnwESscbr8/FF2d+x7+TuXbZP84G+ciFzDqjsojtTHoQTyPnSq7sTSiHiEsjXwJ5by
6sDxYgxOZvrgVoiht2EMhD6kmPz83xacnrhVBDKkqSQdvqrHAqm5T9zQigJicGYoFLnadrw7WJ9v
hIrjTDgJchDtBUlRfd3hWhZwuHIbijKA1XrDpNkQMLXAMZb0MrRrgepAXKDTxZt+rxJnSLBHMoTI
3TrFm9snDVEsIPkZXu8j56tWXRQOaghMFUM4WNSvNOFfMJyqGraIzFU+6qdwwiTpufqj8tw7OBcG
OkgvNnwu41Ifk/bHYuHNdro6zL9wcrwNow/SoeY3GuVFdzufia9k5NTDDfNUcAIfSB3XzAw5V73X
7ZoOulz2k7clQpO1QloKIJJPlCfa7VSn8T6PlfkYJx8jddNAkq4mZyk9fG9MFwprABcASPDN6CQr
O/BItHR29eWJbguMiRN8HWS/GL9dOiGRvLVtZ2XYxt8Q+8HVdRdPBdCiyzp2UnUEaqdhH+efx7jW
7Q5TaMyYpJRLzrf87967BdPpEuJfD1mJ8kFoKEZ78Vm6+IAPPscnyLvDXox7mBdpNO/SvTmg5ZMF
owinl60+oaqpM0XbuG+JRaYwOBj6UCys1zi7iYGtc2bS7N5idSiOOnbWbG8crRAl1VMP6UlxOdmg
1rmXF5gwEKMdHpIDS/3wFPeTH+9LYg7V5L8ohGYEfrhm/zyOKweqZGoaSyA4PK2SOKYpvvBHv5yL
Ka65E6irn+ms04iKMuBx36TsxvNBOK5vKMiwDDc2+/OtDRmHKIeZ2DvWqmmIjIBFoC0UTOcxf+c1
miGslj+GkM9DkQQBZYA0JRaDp8ihzLD3EI+XW3T00m5UnzdwBCwgnWbmlgytgERKIw0CSVlFiSqr
z3pPDPzy5W+f8KjzX8dhJYcYfNs1nGroIx4TlsYmDTqDsMiRNehxztYBQpKPcMvafgvx8rVILIWh
LW8AgdnMbSUvV2qw4cXlW3IjAYGW0+fCZOVHzxg1Tjbb5DUBwBLBxJm58Y6p8uQ/yuEXQcn9nXdI
WgZx/bR+AIz8yld/54l4T3UvNeBe/3ETZ2+ucg4VyJS+4CSIJ+4PHv6Q8KsC1CaJB0bLpLrFZUxZ
Rj3HQOBKfW0sPfsUXDDWBpDRHc+VNgwVtqXZjFkSh2RJmfEktQ2VaRh0WvNFcJURyPtv+6UnI5YK
6Cjhq1NoXFYpWMK/g6ly2WZPVtA6yAGnWXdxvXl+PBQEGrwdZDHGWslqhYOUE15tIglXIKgWMbGa
8yLbovvA1fe5e0XaWFTil+9EELq8qF5Lzdzo9A3IF/gYE3AwxMaUI17gZBMmM+SXkYpunIjKp8G3
ty/IkmKHOqrGKKif/oW8jSQ8FpLQTyvF/ao6WnFKV84Rmh0worU8VZfbYT7/VQ+kebGNx38zuNTb
NqFfEzs9OUH8Nbd9Iqo8bUfDPoJdn+7eiTE0eCJhVKL7M30gkytEug9VFVtXFR8nWI/jPy7To/G/
neiVx56rx6Wlmw2eD2X9J4+zVgXu0rcmUO9H6MLpq/dy2fVgZguJMk8xq99eybmX8L4dBCjBtyzo
1Hky5g+BOpPQWzQs54JKVHQx+IGJgLDMqReVbyykPC6Spnw12cN/0Sj9e3Qk6IZ2g6VoVU4hiK00
rT8T7HqMTPwi9BEpFQ0soeMGal3O73V6m11aoEVb7AAAZU+b+dP45bv1Ayty2fSMayUk7wXg4/iz
lu0/7V7eRLj1egqWQhJcQ81t9E1/kF28ePHQRiAh9dmMgmY77Tv/PHx/WEdqgZwHWzj9yINLRn1C
CVWtEsctuI5qPh+ZOoxVMHRMoy2vwJEWL4pDipIyi1uqXftl8CjbwqduLvaQCqhigREBo9WlI/2B
MKbz6aLVeO6EZGvLirjzeXamM0UBLGm2duj4B6xVxtNY5acBaltZnxuXjFYcop9OyGBIWi7t0ybS
9UVMiQLva2IIdLRXK4jH+QFYh6L9yvf9lACqv0l2xko7pfg/cv6F6x5dxYYt4QFn7dCIPuM+/pOb
Z9YBn7+iIaVZjrV8Aalql6UsNGBeKcKukEdRkDibZzB1Rre6edZcOdt0X4XjE/57V0TtWHJZZadQ
2Xp6IrWXavlu4URWXS+AxTSQgU20YPllRfS2xgLyBr6qIl/uAqiu0nUpPUDREWjZzoNgYyp2gcMV
j/6sb7J977xOsScezfuzzoXjz/1qHGxmPtx1tKOmmre+hvph1EspgaIv6LuKQpCm9QMTflDEFkEd
ajzWBRp7hwwOLYT+XnQ6/UH8IbF4/THuoMtJ638ZxITttvelsfs2HWsWCMz4h5h6ssu+n9kAuKEx
9KeOxUrGGKF39mX6coh/E48l+hdXQZNCTpaGah4ddfPdXHGxMJjcI/28uSA+8UBPDiMz6163vBOK
ajAvkP2hJ51rajNVgG1xtIRNgsmSN62GA8ku1sMCndC+WexX/aBrYsIfZXipKJCk1eFOTEnjlWn+
pOVpUEPmBpHjFs2528ArMRU3m2Sq6cCX+DdbJZW4JFuB9lA1FYGqYr+fiO+S1zSnsELHJBLHDzEP
989/yBdcnhuqBvSo9Vw7wMQ8bNLWOk9Z4gb10uBRnHOHo5U/33VsvgULm47gqQU2/4T95VsA+ZeU
/iHFx2kSy3rbcfiLiOR47AY4x11b8mZSeQU+RaM4NR1q+RAAqGwkJIWiVw4LanMN2yEg9T7Q9xyp
tPJew63MLI+ETRQwsnDixdW+WQz8WHO6EAxlGrRyHkpqu84BDD/t4cIRKh4B+26jYBLWfOWFHSrN
bSo0Qo0ttKSrKsinyDVTFKdv4mkP1EQTQ5tURpx2X4Fv7Ijj53nOGZB9UGsjdd5GiuH+ZKIXctIX
pefBNlyyYm71kjL+swY+r3F2lUsdDvhP+PlawJdwdY6pWmnEn7ekFXGmCZKpesFSxLI2bQr+vu7K
+5Cp9cch7X+ps6PD+qPrTGUkt9czByYQzgqiR7SBbMPJ5vrvnOgGJP3NzcXVyMzuWSFLTWelTeth
PVWFq4VVO6J2SckGnCjWONBqhXRqgvVgHy+2AM+U372zf/7Fildi+kRks7PGHX+bL+o6y+4w59eS
526UL66bfVkVuJLOhjgnCPkbM6ip6KwyCIcLrlw6rFjDzoXo73ECSbYDhdD9FrPIr4lPmRyV43jV
OMjZsOGy+A2oRV3ybiTgRd1y1RGwbfjPqcnm95kzoiIKxVsJQ6scru2oEi4Yb2hw+K9y+ndOWv5v
xTO5S3/cosVnNGM55i840u2Fqh62INeNp04NfHwtN4KiY1fJ1UKcPcKfBGo43mL6eT7Ov3MVpLjE
264gyYNZH30n3x6EA+h9SrmycxKQusBMgtPVEUVPOLihe66ifp28XR1MtVYe5vzCo55vdWxEsiY7
rLss0DDtluWrdiCjSeWyc+B/YJPDLZ32Siw1VgyjF3X1zH9uy2KLCQW5TETTnn0IhEONRCV2Ft4K
oJ9HXyu3ZTQXow8NM4aaJS/2Mj77KKymnm1WFe8GSWdTRGKmKRmgRGv+ZxecYQy98I14+hti3PM5
wgzXas6P+kflp29k40iBIZHUXdgYTYClhrZZAgNjXnJJXuLLEHl6R01tGjs6TRw8mPaoNIkRFGDK
Jk+IRGZ5kIFBEJAuMGaD3txAPZ/eac9y1n0n8fWvdSNSMjhUq5yosroBdtb1GP82O/FBRrQgSJkN
Tx3O7/QzCWdhObt9HkXev1MTFVijIf2yRK1had3j/s4BUDnwMmLj6tov/KY8h8pTpKvcYqYrbPzU
+eUYgk0dP8Ne70xS+QR3OvuLDoPnXJoz111meNpjlNfqFOi6fnLf5bUU9WE/M5pbrnqllzbUwV3z
55nO4C5kH2mtttrlFw1iqrB0hQPzRmagosNonbtX03frm+lX2gQXxNl4sAI+G0Syebc1KLzKllD8
QKWPWGVkKr3xpGKT7xtliSsugx+4km9OgfZocX0KcHUxC4N2ql/f3rioMB6/EELJ1rW0ZYFQqI4F
rYnk8NdIagPj2KGZmZoHSobaS/2asVl5q912PlzAgzU8WmyyZixgNt6BHbErHrHh94qL6cd1guDL
Sfl2dGRWVhr2exMfE+yDtwbsFnBMVbarA8zrCaljDglK5ItYkK01L1RELs1XmCORrPfXDCYlQuP9
XT9uhtp9GRVwchvSs49qVwueBQoLnm+8JSNeXfR5878zICE8ywWnntj0XTQJTnmCskEbbnlBuLy0
kczjDRec3FZS6abGuef7benOtGlAukiqXvoX2KCqKey1SOmpyvXsDayJYQdyga+ZjxbM0m4qJYG5
3jY7NvfYLRN99hlpiJPSdsraJ1KeSj+fDlMGOOTjt6Qgye99dL1wKM5ji1ysFWG0cSU95vf5cC/q
v87UcmAeHbbCBww9c5rrznIJREAhgBTBIm8yLfsbIwRm4a2zIysIuCrv17PkZhC+SFKwKCV+GCom
dryREZxJMjaCIz4KxkFDTU3gSTFLD4YadJ4eacpJPA6iewxUXtOkRfa59iS+RFavGKKN3JSbKwIS
CdeoOfLjYfr2rg5MnYzheB/tXaUURUZeGGhVWVzEQWbMMmbNYl2ivRpl2QNvgP6F34dkJyv6/4oM
DbVoVBFZwFAkVZruLAIAc/d56NQzAlAD7VQcly8KlxKJ4UDiE6Zf60/4SCaW1JwAwdoJ8PAAZEx2
D/3fKpGU+8x661tNnN4+ShpsdFFrjicaeO39Ac2JHuKIeOK5pi+KFk4doiUiN32nl/OoroPVwIZL
f5fKdFa/D5JkFTD4z3golqWjvC5OtuBRLygqy4wuds62S1VDJv28uiTlrcRbq/mNy/Ua/EPuA75o
b7mje4oMZGHX/qlvDuMxgPzR1VeaazF3Xz5V+ZswTWv0fJSI4b79XVf/+D9EwIggIsO7bdJDC5jt
izZHGquiTf9FQKuPzVsosrlC6i6S9KoIr7tOSc0Vi3BcGUbUKI/TILSv1fTKDevlLtjDp5yu1XSQ
qENNyHjAQDQHS1jeDUSAZOtZPeVJY4EEEzKpY9CHXxU8uAxT7b85wxcmMh8Uhc/RUnf990zA1Xih
pIbVHG5UXMu4hIf7XryhA8DKgGwLpVgW+tgx+f2jEUFiEM5lN8ZBDCXV/2OBR7Jktm7MnmQoc/6a
kUNhF2M9QqQjY2ipG4g+jtJBffm6cuhbSTvRScJs/x6ccqi+poH8gP8/x+5heFRBDN9L2QQWkFrh
moOehmmT2Iqdi5Si7+y+niASv0HumQT4FwQjSW27ASz4/m9eYhYN3ROv5eVQFb8sonzY7XAIO7xZ
i7zmnnO30zY+DZK6PlgsmrxHluW02F76OX89VtwhmU0e4gGFqJByWIy1t5kYXE6Z6MFBKv4VGeWy
E3kUDd94I58QsNPGcH8W/yNlqbg/s5XSuPUTWwbft8CdKamMviGhWgYmX11ARqACChMYeoTNyZlI
YainJDQEyLEP1+gA9IuxmwzgtccsUHyE4H8kamItyWuJnZ1e2VbFoo25jUYY38u6U3eA+rDNQRsV
C93cc6WriHkR7x70/fH9fNzXuFpD3pUXu0EUNB3nN8VPyLkIUJh+JKnhFiTRPPvXDGaHnThFlDmn
/RgVmGxEIxctXS6fufwsmXWk+pRkTpxxYGv8MMteGDhOmouv/AKLr5WSTpyRTdX7jPumDmIUEQAy
WTMBkEGBsL1c1VNex5J5e0HtiF3aOAhonZ/ZZBFBw57TTZm3/LOvdaXVqrRKkKFofAe4ohbNksYG
wn9zatQCspVL6ARdPfiAnRWGe4ZkZvrU2LM/Ak6qAaWt6mvp89vZWPho/tAINijskILuFDiJSPm5
dO6Y79+WjMcQTboQhRa3JEq3ZqHLpl2lezG/gbS7pjeLPmRH6KMyN3VFGWkVB1BWDM4tm9xxVde8
etZ1q6MxSvuCu20FLuN9ouvWsgk4mqsiIjEodJ3OJ1Wi0BAnacLA34D4B4POI8ywCRY2NUqPJDa/
uhXJ3hM7kqQ9BrICoEfjbRTHSaT56eIvmQldLjmeUbnl77htpSxZpnvsCO1W/9wRHjkPsQi5HLAq
7owpZ7nT+YnzQZ+uc8YzqdAQ+bX3Rarf4KHuyolm+bdWksNOAC+//pawC84mVOx/B/wUwhLlB/4y
U2J+758EYL4o2XG2qTGH7k0WbEwgHV3JcC/QrJw2CsxnYf+Rtc5gSZOE5eT1Lp9uIKRvJPjwW1u8
TLJHk0DiqTrobzADkHgSFUTUlPyyAHpPlEnLE+hcvS8r/Qqg4CgKeVlMEFe8R+snsoS3ZG6o05So
HEidENRXLJZGNRhoWCGtpnn7Gn1QHWJ/3YsZehqjunPl133R8rbIFeaoqV4/hBSqASxhYE3A2MSy
hpn9Ngt/P8NEo4lVOZ6iIoKOSZMAACvQH55/L/xF975BxYCKO9T8+Iaps9y/zqP9jeWRZ70fUnW7
jJsSWImPgohKVa9wJvez9j6OA5OziYusRlZG7qO/X12vcVtPTS57tQLwOtvmRvPHgOBct5Kxdg9w
gycw6VCiWzh/xv6W2xlW0KLCj+4LMQfSYVQC0AdLb9iGsG6qVjxXkAOVml0q46dawpxvchnBMFg7
4zV5c6O3VcBdgxQIvEPJjGPbiuNu092momM9nlpDwy4Fo/shEqwrkzPVvGP12K1ZDPLDaCbmkAiL
RjRfGJ4JHVc9eAZFJsCY+DZkyU94R/wdm6Zo9Fgi4XTWOkiDKwCN3q+n/fX4sUmkb0o3G2LXt1dY
+C+IcEIqDvC00CfTGCJFJwrB1u5BWvE2O3b/Wg+J+YrEUzjRd6GCuaVd1Z2eUMFhy7AN7jkL4+MK
LUe9dQcwNIsc3T20kA0kfpLo2ZRgwRdpgqT0hB4w0U+yXCFPEj8pXVCpkgAlIxg++YoVaGQmYj9/
ivuwYIq7y5/vn8thA9tuexl4P9SLY/4f75VmaFBTU8UNm/UHOTXaS3XtwCNPoPUUMlgyJyDdZJFi
IlHZAjSLi4QjdrrqiDXDsfsPLXOT+/kz7z8Euo7ji1JVS+WEy9aLw6r+4y0A+uJ+ZT8d37HWU0iJ
/V0vZh8gHST+NIJ9MH0oXqs0MuSyZynWZOBrSPFAFOfLjAImWM4VdiaPJxGNuQJA/x8DzDFUxeu1
E1w9VrOhKJbP9d7T/cE+U76OCVWTZD3nxTccyhfj9toswbZbWfiFDcyWkG/mvzeOJoQP90jeeHoT
NbbH5BkIoMaaZ9PskfCIkdJ7ktamtPk96pWp3DFvzG691+fwLGZIGvLTtclP8IDWXn47Qnisyp51
HjS3IPzU9Grtg0pbqe7oZDAV5OE9FI5Kblg1BDNaAI98O1eJbVyI3BDun4MLv1W83ChkVYIhgp+R
P2MfNEsfn2Yplm6FwYrY65gsbiwAyNC2LLexnxDTTHE560kO8LFKstLu+7nkYqDw88ZYUXt1dmYP
O2EMmjmN04Cf36oGaqFFVUzMcITnnVg1SWRp6BmqaDxKzo68f0qnJx1XrOkm8kMkRTyvMMgMRz0X
WbeDFK2Rid2lIZW6gXgJ4zJUcyBFFwf75I177NQyIrXSPI5RblIsnkuDADd+JOnydhPPracwbEWF
k7H36vtl/zpJGlpeVYj39FLlPHzP7lEpznn2fsFvxceDoIPKyL8EtghkSdTfZRaROLcRtAduYqdG
T0qpy2+WlZxOdO4vf/nyYJKboNAa37l6JJ5uQuGdMbinL+1v7t4mlHnVsmprKV6S+xIsCGx3QIJa
DhucNqUMBLavcEdVkNlajm6Irv/QPlbo6HTZNv/8YutWGagV3ShXMk8aPr/qmPFXaLaXNOZTb6eZ
8xS6SBeU6hFT/hw+mkr3jEpEjMbxTwVqk3Xg4H+ey2H6KM4P+sxX0yU+XLaHT/lrtSn3LoJ4KO1I
3NPVJ+dCqL7j5/cMgQR2d97PPisMfDKdDWzucGSrfZsIXIUOr6R4NT6Y4C7Edgu5x4Pnn+odhLuU
4v8+rwq1wuFdf2aUACmyGse4lVCI011HaY5wSsJOr3p/909yrzNEiidJsyXSZCBKG/NbM4xUbFj8
SYkLMi4k+L8BMQ8FFXkJqIrmAbOk7vemMYmN524bMjz+Q6zoE5LPgSTU27203MlsgR3vHaIuWpNA
PBPHMVe4JZezMmqDw0ilCsa/QjIE9j2w/HCttWSVwLwsRpa1gBDLho2bEpiOIpdA3OHlsA3YiEA2
nBJj+0GJPiSVlzfCkPfWj+ZyTOeZ3L3SvHoObP1g5Er19LZLrWzkyu+aojUcEaUJBjZG+cMcuubF
Xhobje/4sVfRVEHKcw0lV4G6RQrpGJmTvFLYV7K4uKwL2zeMI0VEVTq9ZUeAAU+mKLG45JW8DlvF
Nd30cuIWmcACtTMpves7VQAkRJvJLsI+pHtzzv+djZDS+UsC5+zIHeKdx2yk/GnKFa/XwHdPmm/t
sBD3i4MfFSXdMiKOXxBY0YqHqee1YPuvt1dSgbsJTYbF67dRXvBiYOegWXJuOW1wnwPTt6Rrm+bg
t7uMjRYSAGPIxgyHfTKOBieooLTQJNZiMkcdy6+NW3i4ZfC+CVpmUM8pl5UCVt7+1CrNwU8LLuf5
qPc0Ko76xysAw9ft9o7nnmdSYUXNWZHH7e3P75g0WJADKyo24UvyXOIqWDsWPHtsyaDdcHBljn3u
w0zi2H89S3oG9EKc8+qSKdG/v4VzZWKkxx5xiFIs2RXqyPs9RMIQIATcHOUoAJYgDhtkpQmN6zB2
4BAgOprX9NQG+xQ5zeOl9TSXy1TinFOAHAxn8iea6dcrQZFUqG2zYfiwWd5DfWN/BB067FleJy/E
4d2JKG4cIv8RM845JY3Bi4yLPvWGbI/4AzhPf/H/gAjx1M0FRYUfiJfcpLWwILfwgHauiH8XMZZx
Tx68Nhs5Pc+IpwtOedd7LFPp0nATlJFKcYlaI1zBN3VFnoAbLXHCrWRtTkx8pxtYmPIgGMYT7CDk
nDcFkYhiJfg235IS4M+/T2Xwn3Q7WUWQ+l1iqJXP8AFjG1HxZBCnGaL1D/ZNj7y+X2vt7ZuHh4E0
9qJgFP8yGHvfhd+DONWsIufw+AM0u2zvpcUEzFm7/373DCBl/DXdl68FIu7LNQhy3imxs6hOxjcB
fMxQI9XNlqnR9tVqkObzhgnWGjTUWvE9/FIu4AiN/fv8mgz5QGqJQBxJvCqK8w51JhQ5i8zrPhWM
r/YFd0ZddUFsX1/LNAbE/3bx5CYzUCMx+sGyGw0MjxjGW0CsNeOGUxs7JshGkYw0cmC4lA+RACrV
19eHDPwC55Ag6bNZh5Cq/VgSMDOxYgjoh9laiThUKqKHXWTvrPdbuO20+RtSLsQBZGt7RL0qdeuF
Fvg/iFDB0xsq+5T+gWCmracUBWfXu96xrDQ8wDscuymwHibihDV3BKrRhulE3o7NeRuCFBXYV6ep
XtYMdtQ+CnRK9nVSqMCa+yNGfgyPpS/+whUSMySO3wXwPaE3F1lWjPg5vDUrKPnYOvAlCq38qrym
5rtV69FPEGJnlfy6smZ9uvvmRJkuAhywWwTL+j5yumJoJSQL4nDhn04/pzK1f/UnD98lK16mFwXX
FL/bLT24pwcoihuyEJB3aDyswF76FhiTdBqVI1iOznZv6KdTQZrjIaaJZ9RvrEvaOYu+7w6fRxx4
D3VGT7vxzw8jWtLHJujR5KLM+M396jXfkb6osTZy+RY7xQHa5w2O7xuG3VHZdVn/EOb5YeL/RORF
dfaa7t6LTfKwvu8I9+OvGpnHTbOVeIu0/ml3UyYBIwq9fNc0vXZ2Kr8lfRsUXRXtLP/BHbYp8P+w
vIQ6mh8Z0uck5yLZxbFqYN8cYa8w8/QD/k8SlB0ZkAyMnW7cTgjasU4K54z44qqXC93qikjOfbT+
CW51WqH3yDVGj1ibmz2eZ4MsbR7dVxjJF1cIJdChjyOYwL/xeY1LaLuD6OzoJRg8gSurVaI2f6Q1
HSjCmusTU+dvluXViNdEdFVYbzQ5J5REI0344ULx/j1JDos0PNT98cwngNuw1TlBklLBsV2OzCE8
DhWeIL8r/cryqgZKZica8fl+/jM1Z2iqufKZue98Y4KTWb4TFtVwYLQbOhPf50ogeGHJGA1ETQu6
pPrBDXBMi82nY6iK/pHOu9VYO6frKPPBc6w+0emKen8GXQHPuJaxMWC0j8dBAY5/FyGROfB6rYps
P6EqvyKg4Plg/LCXWhAoi4Uc6KQ0BLPIwCFv33TpDUM3HxOMYntPEYJHiVB1DweUM4zX1Ov5fYmZ
SqHWSUnPnzwvp1ZfdXEAg+gIUy09OrLNylPNvvR/rb7X5VDNvAjM3dTb73uyB0sbCBljSMNe21V0
juxE8WIb7kFd/dbXCrVeZJl2oFS1CxIS2Eg2sTYvjBg+Oa5NmnXyB37K86TC1rpugayhW68OwsVO
M8IYwA+nYCqmXLHYppExx79F8ZfIPcouM54YRlz/Z0NHtt93VXsP07u9aWoesFlsJfYaJitHMh/d
9AUzmLcuRrSq3xL4u0RoY3hid/BAAD/HJgrQH3nFxsJ7wv13jWyFHXFbcWuT8DQ73vPycSjsYn//
xa0IQdv1RHO92DT3ctQyVLukhNIo3MZ09zDNwaJWaPfA7CBv1mZWjUNhAMzrh3bBokxSi5e/7J05
5uEIiEbzimxR1w6WAViLvhkZthKJHYcjUPT0uf9h1mqs5LFS30p5BAh6C6jx/j8RvaQMBaVHSc7V
srBVKUHXo+++U5q0XPNSaRXvslHw0vRhNaVjZh+iQDX10pyEqJqR3gJ9CE6YxTfVkq+8wGtg0Uwk
28WOPrczbZh5XS1NIXcgXF+14sOAr2dPr1QxUYGNY+OiM5HtxTMGtKDUzTAJJVukcK1c1ZknCwB3
QpGgS6AFiIiR3nS/jK1y7taBnJ6FgkLn+wbMMr/fYwMtFAqSC8ZpqMHeuTNZbOj1a0rR5g0hkMOj
DEKRrJlnzypG8xlh0p6lcxKceShVS9iIKpTDyTse7iYidSXSjcQaqLn4/DyF4jtvQm/ZYjOgbGLU
h1PuwEIXPsP7LrNeEr/UPDW4e6RtPw+xDJUHGLoy0Uw3odNMqa1nWd3XKjDoN8EaJyMJSdPdei7p
wN730OgY4MQx2BG2nXmPrySDpsaHvcVD1dE1rJ6jpYQGXNO1hsppsJ4abCKLyed7PkZAYcyx3nEk
L6E+9fisBtLq+p7f45mzOSICWlDEgyTM092IgHBpQI5mg6tDWyz+KFmIQl40m5jYuthsIKuvtV1J
tYZI42K8+hhE161+J1+g8VxGU8h+E8yjE0ORdKriVv7+SEkfb2i542sUgsI2+tmQeIZAnidndbv5
DLfzl1s4iWtmjtXUxGtYULoCRvdiyyQuMdIbUMxlpd1edAVK2CjrF/LtY0F1cg29NQWNN54IRCTT
AEahQ4vivQolNQwq+hrlMMNXUb8Pqh1AdsVqsE2+F1a6ICfakSnOs8Xt4SQ0SK3ywHMnMFfLeY4i
To+9JD6g5Gm3rp7KqRHYt7DaJBsJVK5ls+PlACLfgmn1ADnvMmrt+465SEtz9YHjY8TKE4H1zMdZ
zuNyB/1kuQh3TwGynl8Pn1s5COnQlcDNrq6WXznJ7/1XwWT1f2R3ZACFJEOcGBN4G+k2ZtvH7AwE
2GYUM+r2Ky2/sxQj6H6hFuaN8ToqzLOr+5NI4DrlgUfIO1O+IaDQFtcavmGiWsHy9pBaGOCgjxWK
BXheEmKKie/LGTuv0FSFmIHL9cfz1pNQOHqqP+m0D8IecVuvgubSrQ6KRKOEmFFGbqGqoWd5Xh+b
7nykJd0fvs+iT+zL1JsBz8MisCucSlyiZrZanLeL+5XcRcCY5gYEWDLX+19LbOCj1UELUm5DXQsi
504PPAMs36h/fg1/zW3rE2b2SKJY0ITpTnZYVDqxUMRlTYnqstmEY5/yZvQi2vsRMo8ulOWDxQRq
8Sxw3wwLJxjvPjuWh+1mQ2n9Mysm41N6JZ8eUgMd+0yDT+1WFSDiFEZjjpf5O7yN+4fW7DstR8P7
swFBO7NFXwCvAcwKKLBf4Lqb9sJ8qxxPmpxyX+6IWmwspiEL3/gTn+f3WQyOWXU/YEODJqtOCFmS
yOnuh/qj5Ob5lWBTjxD0jQB/xP83S7PMgutD0751xDNls8Bq7s/D5p2FCVkuLfKJEI1iIPcSwMLm
5V6NlF+OVWkjmm7aruVRJF1yCOJmKc2f0JAlIgRz8yEu9+DJUhZ+dY99kJzmRJQjQTxDrg5zdPMD
z/k39d/7gMefyDZULZwcvJ55tuV9W6nx9pMsH7BizQ3P7opLEsOR91TvpVGC6jRS0xd98WZe8S+Q
JUNHIEkZ4Z7HZnO7Iibk/ww9rnFnBItTRifJTQDZxa9kdvJgKEPfClhWo+Ay8HWvItVlrmbD+WT9
oCTsxttYxlG63kvA/LkPtYsrhRwFLXWodGLfrLrSHHNP1zM2h/WuzBz+XrygbbgaZtRFw9eGpjvU
IoEchuavfXcU4wHTEwVdZyIUvYecb5QJ3dBgBFIz6hTyUGKRs2b9Zc2Nb/dvL4dxroyDMrJ0mUR0
we9mAXd6LKBDkzXKEX0QQVpiPKYGN3OCoEuWqZmXuSeFFx+CJn3VXemI3wgaSk7UnfShQspBrfqM
8fpN0g9HOrPj69dLy7LgYbis7Ggtht8pG52eV5fp+OSQidTeI5Ri9cZl9LMTd3OoNETlMl4ERROp
ohGZE5cQE8zbTABJpAFmMnbLs6H36HavUBS2Fn1r9plDrbA7IC4W8mlLhMWEYk3sZYEYTBLPtjzQ
yPROhH+Mr3jJ4aCTzwLxo63SqQfl+ZMMcZNEj+g+qqLm6E25Yed4ya6i8vBHMYUxX4zQTI7Hd2rF
DQ5sJRLR+rho3v2koIqHcZMauyb8RLCkppnATUeObSz87gOe8IRmr65WY/XkC3w8dMPF/nWeUFtj
9psXOWNXT3p1FMYH+vRkWYf5wxszUPkWOJmLPZVL1Vey8iYitpTLV3FqeTB/tOC7E1IIZMxXNQ2n
WWV2emK7s8wK/77IJBhmpAVlpEWVuDFE1GPWf4HbOjqsorlw9/HWOqKb2L3JTpWDgd9n1rcxtWIA
dP661W530gD9oRBAd42WcK6KLAjUgj1XaGfQAO4Hbrmf6y+Dix4HSzp8cAu2wBzMt3Kp/95/Mb+9
5f51JIbaSlvXnG05LL5m70NbXb8TQrLeo80o9PrCt+XM1g9A2ZxUD4W86fOKpML/UzFfiQEz1Xs6
hC2d6jGH60NscbEv62kOLlb+FHXa4Kv0gNPlOsm7CYrNxie5XfMxNlGsOSRzkpZ8a7fyzziUIFN7
SakzLKKrTu+DXXxHxwI2rH6cvB2pxyQ9LW4mlLIPOOJZe90jobDBciqRQSSPJC7za2mODRySEa6s
FckAuqx/GgOdrAiLpJxCJL/y6VrzjCCpjXvdaBc6w3du4EBr4+sUVgrXAk3SzWHt47MzTViUVpWJ
epbWF0Ivd+i6fTooguyWz7FosyG9WeJ0qW4fxH4pZiaCdEVRJFtuIvcUgQRZWDglwSS38EA1ISKg
lxDreRnRlFS7i0YuJspRQRpz+79+1DiAhuGuwIJb506p5yv4nZP/DoBxL9DyqqVm7VMdT71XJiI5
g9XT4MDMDPiQb8Xv4r07pdNokSolZ3PB5SGUnRB7WLLGbgo9txgx7fLOTPxlltzgv6ewLaCjUbzE
lPe46qwDhxrKmCd/cpagUJbNR1Sqdx0H4Liq0x0wnb1zJoIkCyZk9P5x6SiIoDN1r+qj0lvr109U
z7QDzo67/CloBG08PR/s88o+f4Q2CQkALZxVtvGHY9tdIZUOAH13nKzUOy8kkPmQUS1Jpmw+eOoE
edVeqhLHz3Sq4cFmSKoTltCAaKHEQbmq+lX+NRlRIrtuufjbrRcpWf1EPKSlx9FyxJyO91FNUaer
v+TiWPG/pqwswochZybhQK7FQqTMAt/ulDPoZ2JTFDedgaJhSwcGDvYqf8z1qkxtgjCy2YwOpQE9
zrwHHTMNJe1WElQLxcJPmPPk1ZDoCV18Hj0egrDllo4PqTX0thIHVlUnqnW8DZq3bTi11lh27Xdy
dtT67McXM0xX5s6D2dzxTLxlEePCgxKPOLU18+TnNqP6CbVGEo801c4HPJ7gSu9HVMgLeNcJt5mF
fyN6+FVuPldz7yxOEv8oNtY9gMxkTLTWWZqP4UXiWmVPuI5JsQexX7XGoZtjbJoEQQxn7/RhVWki
uPAUcDz9rbXJLo+MZ5nUXFJqwhQ1/a+VO8o616Y5s9BupV8y8FvUkRJLamtsLjvUKVKxLPwarpKU
T4Wg26CIS4kY3vxa0KadNjKxBj7RwM6bufwkvswAe37jiA7vF/ROvPy068Y4Al0iODrR7Vx0aVBX
fqdFInZezC6E31uQ8yY10Eq2oGfa5Rr7T+vaijjvtmWYG6n5eBzDYCkrnSPN6WhqoZr4j6QmG4AM
rE4jCAFyI00kntWq4hTT6sDEiP4W9UWLdVUI5wnHlAHDaVjhvnNtZIrf7KPVbenSDzsAlQOFhK5Y
6X43eZWOasW47Ba6wSwGpAg9Fn9HuzRvqiMUfjviOBxptIjEXNXhAtKtPuql9NWxS0BJt8IzGNSv
3bzL9IIH4yJXzj6isY0sndcle3m6d9PUVreWXEgtqrt8zhKJy28b2L5V1LHy83wSOU5UFLvJ+FP7
o55dkC7j/X5k21L/H2LGsHVI4sH0oKb4hgVQSCZB+CUwZJKvfnduuC4vKMo0Pe+/SuOwe9apxgdC
zi9kqHcCujXhhPITPOHARhKfmOzidFxXHeWB0FIDIPbyQMmZr6O2wga4uGltV3kJ+JfRQ953Laon
lbet0Fb4IaM3+/gwtJkfwzzVizWkqxLIIkLYHtxzAF0cRe/LDmTMmHJj2R7/GMI3vi3Bj1TN/IXE
vn04LUmgeqxSQbIH8dYvnprdbKjAc/IfDexGsO4+Vt1ydd1F97gG4vczTo37y+q+iOuJn/1tqZdO
1LSBLaHvks4DR7fRZvr49FfPxWxmPfXMWpt+J1G6Wt57T9WT9S5f41vtfs26vsBRp6/Sb7sZCqBZ
injGuPuPPNwf+w1zdzAK3BR8TcJpmbenB1iahkxjKBGmhZxSczO0wicCg1Vl61cEdl7b/U4TV8g3
Z6y9a1lHpLPfYR+j4y8Wao8BijC96AQbgnu1twWD9ylc+AHb7nRrdGioHCVQDzrKRc8FNA3AwqSQ
YEDkA5yhJ1YN9HtcDDgnrlsLgM5HpPP+vd1jO2Zw1q+GQyS0VIHEPUa9srn/0tYV2qF9bH+ldzEi
aJNetkHG606DIuic72bciwsgVOnjEzZYoKq4i9Iqg6RsPMF9PqUHFI4V5dQ8Qy5LY0PyTIt4wgnv
ELUMMSvlWeP7keWSqFxAx3THbwxPFj1H8ml2Pj/7xIJhI1Sufb9Sgr9lEzjWxJj1MiTUhNe7bT9O
J7Mvp/lg5yc5byiEgskbvyLBX03AFGl7UGTjC5DIxiwR7AiBM0QJ0uwCQXYgzeiXhXJ50XUSXjhe
cPs+gvcX5+y/YvvUyz4dM10QJ9Wbyn435+EK2D8cSR3j/v7AI1QDfRwaYzNPRk/McSHT6+4uhvaC
2MMvrNPQ5mUbeYknCRqxIfDZYb0JzG7tTEKmgBhKR4KH2pA0pXlbzTI8zOJ7FmtkHUJyetmwQA7m
y2P85olAQm/vhF2jH3OK8JVcFMN6dakLeYHkQjrFBO2YGNLwbfxjXWVyCV/M4h8uDagE++qHZCEv
vGIEUlUYw1/KA7xoxjwMsZvXM4x84VHnHa4vGU638Xfu9UBBFXmwA937xxA1JXLrk02F6KYMPzTB
YNlBJnWyNOpx1Z8857i3bb6ImvTu/zCKQ0N7vSUp321qfeOvN4tSsYN0lCXrOEdFBPwvXyzJrm6k
zLt2XKFxf7GKEWJoQD8qQg+HHjqzBoOsnOPgtEuJHJ6i7lp3LBNuiSux6ulZwegAag4oWq3PIGMC
p3wl+oMHMkWHRKa0gIhCLjauc/UJN3pb8vXRoBciPIxeXD39cwkE9tvms/IeEVbgUNQ+SJgJpKQh
YunDBmnTzklJxiGpFTkGjxLU6cPV8rPSLzSKBq51htKhdFOwwv3aieM+uJ8J0LfWglfq9XT1xARX
iOrZSGsQTce1huqtl/yNAGwfB7t+AMHv1rsNPTbmaHi8tXcunZcKhImIdxqhrya+NzEvMSOmx0cA
BmSCzyjUEC1MwrbY5cFB2jXAZY/w+acvlwuLK1UoF2NgaPzL4SgeNX6JmwKMp2N76NVPmkRCF2dK
QzRgegvlNkusjVca4oVIMZji6duUAd+9qG874RubqEEVlcUWWVLplP8CaWSYwgtHB6OlrUEQjXjR
yrO58/R8gabUAuw3AcT6ZWce0w85Lsl/j4myvJrVL1P36xH8+NLWWniYUVthtl/ii24Ssunp+rEn
k9Ei3TA+oMlZOhyyspgCmctYPJC9IRblpGNY+92aGgZUtEjgY3uzUc8k+GMyhx4bywJs8+9XlxEe
tjaSGprggSTjJSJOA5i1ZA64gP8jrH/L3fNmB8QBlZEBm/DtfpjppcTRetBcceUz0sDmO3Gl4jO3
pxolumOh6SJufcDkEbRlMbxVVQmG9tDbQ1IQlBNjS3SHZyXgNa2AdxPjs/7CsstNNaezUVAQPCkp
g/nzb+xAHQ/xZ/ZWMdh8bz01NH0M6hOWiKl5s6cpHpuUHelRrjypdylSPySzGqMUS5Laob1nZ7vF
PfHuKgmc6lHj5llO/JdLVpwC/UN0rIVoVffKX+My6Bk1Q14HDRG8lu4iB7avipjYGvJfUUAYDbHn
9SnfIca8DihaubcYk+tXMJIuAus7+nQk1hN4UjSj8ihcmmvXuA9EDlViC3RiN+XwOXBEbtF0guRI
qUDdNh4EeA0ST5dCIAYOqvACkznytmVazPNdboNzpyn+AcF7kJyvpvFtrwuErA173Go/2pdOzlsG
8wyL6dsT7B5oeHbbq1NvQOZwGQKs7g87DVG1DFsGPI2lA1B9m/0s61dRw8LxhVb44NSK/LLZaObM
oCldH1nFdLa9J5TanImGMDrFJdA8uznBVoxcCNtiVZQTepbLiw8hvbjC3kyDFd6HKMDYZMK22cZJ
j3YTMGLu7gE2YM8jzVcslSV7De6ufbrhwLEMoMugFx67GBkK7EWY23PoMQYrbbvEyNJlFHxhOcX0
5/s/JhHmrJJeLVLh44HSr7g/x1cu7j9Ze+5zxjnOsXyHvPGcrLIpp9kEsss9/lGXTitELritL6jk
ph1b2fqg3+PcFjDh2utIidbS+zDlj79jPHd9yUPrdjTRzivLHvh9ZEKX2E8FjjE+rK+J6O7eSzOi
ZvFOLBNBvf2PQwp4r2+fnkMrZK+UJSMac9PMFo8Lp3gyK/3TwdbsqzPe4LoYytg8106HrSg4ImZq
Fxm1TfmcxGWhQQGhw/F4HEs5a5dKvC6InpELmFuaAx+WEuStqmnyVupRLv3nZly+12nxxS2vb756
H2DBFuUBAvJfRwlBxvfMJIoqG+JkwUkMIizIZWE/1wX5QUI6lAJJQ5mSqctvmpmZClB8NFIe9fir
TfZuYFyi3ESAFuxIvil0IKgB0j7291xuwdVKJGcBpXOYyzart1qi0hR27u0j70kRDQF47aJhLL0+
EWSTwLhfba18ZDFI3Tjfb6No8LX2pQGQge8mHKvNgR+GucVvxqtjwAQrzYk2HyDC+x6tvz1XODWa
DIpmSuk1RXBmN8UiBe9tXxnOY249G2hqsPzrRfjR1j1ZqcCwSxm6prxm/SkXXSMeUuOWY5Z51Xki
iaaPNdp6cyd3K0ADNba82SAQ4ueTXN4LaqmlB/a/SchCZn+wyzjy/zm5HXd8Dkq4io6v02IcrcYm
TV28L/9sRM6Lj29Qr9aKUPrkh4JqeLgWVDbm68i8OFjOlzankONLEp556tp3le5LIho4uKtOJLFt
sGWFuRq2gEJ91pUhYlA1emqOA6kfX1+Rf550R/NpxkqBNq80AFio7z58tUSf/85TMhH0tU5Ly+aI
g26kkqHmGXjxFqbYJRhAVmRpX7q6L6FgB+rmDe+Ta2liAX1Icmy/pK4Ovx28PvT4VMy4RowytfTg
H9lAvkkXZVjP1m11dapJX2K21z1+bRaq9D0N6LEVi7rChBQUX5ZAqOhN+MwxTqlbPXd+Yc6LTZpo
CQV8M1CTIxOaN1a8wuuj/o2f7/QQbkuIZ6A30iCEhkvVfEAOQq7EnqM5Bjf6SAXr8gAoK7tXGDqq
SQjBG0CRdS/qmI3O6H+rm8AQEMsbXkBMqrZoeE4rbagwmjl7LNOVRK8WkjDn+V4xmQbZDXMRKPu6
kkX0rCVY2UPpCeHF4YgtCnLHPhJxhAvVvDafA6yqJhAN2a+eb7ONKSwdUbNcfqOChSkbtuEzwG+j
zL+D8Dd30ZVT3mIkzp6K+DAs4Tl2AdlnqaurdWN1DY9TiF6pF8pHPiCI4Ykx12eTPKezKwLm1T6W
/uZNqZ5uLMZbHi3DMeb9nNOSrDLWNHciNW6TriJfVUaEdaYUGaK0EJdC836dOpgBtLV7XsIRxChD
oyjH5u1DdYKRA0+Fkj7gVj23k0JXz/uYLWyfyPjMbpb/ABSH216dZbbGLEufSz02OLrsQT/5++MC
UPTvMac3R5jttIg9DnXIjZhV70XFKgXb3EOk+S989B1BMnvrXJB2N3fsYwTibxWRrjJ31m6LNDos
CXH4H1aFRsDwzr17P7EJ2hoWw3PucoYdOcUY7eymTVtJGYZrUkALPeUyAhGbPoKfEQ7yF6TG0pEM
LxFfi6UxPDQn+y40sR4RJUIPbw0yhdvr0lmLGuyf9bsR1hA2R8IgTGtnb5dbZrqQ9bCmm2j7Dua2
7LBlr5Rd8MckqPtca8+vrX2rTxg/PA0JzYiNc0QkmuGTglCw+uakor3ovJ0XdEoCFuTHJy2bNYiy
I41diH64IBt2sWB9xQdPZtvyrL6nhRr+VX/xDHGs3AsOrse0IF+GYiRuwP1sOmqt4oszGAQh3v1q
caky8ev/Qn99azWGTBEXGZBlpZfBmG/BKKmXYaKyHhrFOXxSnnoj62R67+89iAfXwu2gMDvPHz48
5afQjkydNYpL4uZUVr88zZk50u/R4bUPAF2nbJ4xlcU1kFOv0h+QZbhFtbb5N3zTjbozMVvcv5DS
p1QRhahtSGcCYsyGPFRLUXQsb3MeZ+13d0IhHy3rh6kU0WgYZqFHPQdQ3BjeJwQ75os6BG9QX4Au
D9enwOzId6F4pECI6KZjH9sblgeEviNtfdBqxMr2xYj8x+TnY5USZkr3aJGv7oj/quEie0xUZR3D
63Qgy3INCGytAoTWpicLIc1lAy37+xhMeOaZ2OgDOSLWpbfncRFaGRbIrFLe18Dq2oFVvRq0L9W5
VajnQBWX5LZSXSDxOEEpv2F+kCmbK7K/UfWMDWm42UapFN12aFnxEWxueCk6Sq2tdfdQtNVojQOj
87Y3m75Ajbr9e7YpYWqfCYR2qwowEZ4gm7A0zwOduKRoMcMthBNciec/bjNB3A969aog/2t0nrfo
RFYoXA7zm17ZEp7+UAmfprqPutjrgOZooB70iIKRjPaJuepv7VmK7Z1jnYPYRJbcUGcpg+eSN2pH
0aBo/RXTIgW0UTQa5BWT0tSALQCWE+ozgm3PtLWcSeIcCDcbI3T4Cybo7z8rPFiEURMwF7opYyXu
rzxUAVHxx/FQuaVlmNPCOSFD8KjZQ/3BGFZ0WPEMhPIsNKcypD16nf8WglDi/Ffz885V2aVbtUzP
BsSPL4exsf6IPhsEwI5GLIbARLIjFQYRGLg/N8RZ5qm8Q1MjJBPUgRnKGq55sQL0n1W8MVmeZeJy
2MfltlX/2cXIA5vt/liUNrZADAQBBr9NT4dkQ1jluyPl9RyEqg8+7rLVFNvRHJbLtx6V0vBXjik+
0wB8c6BsXiGrbkXrBv7CaOxqCxlKybO0tFHbu/q1Ld820LMOmlgXmSeLe3iJKHBcvMmLzASmOMzg
jimZgLif4ckjHBmGPwY4G83ovkqO4lkYp3iG0oXewnVlGk2phfTSYspdn/53lTpJo/ensjQ0BPr9
Ku4SFDJxIdiglEmh4xhaxS9uDyaPgCWInHGR0XvHHss9HfEOysJB6jT1X1N8XSl0cFpldrI9Iker
ToKlgI8//OmnHh8wy/UhwFGX4A5iKmmCm9Hl/xltBE9yn7z39tsA33KZf4wgbF7tHDZ3I+psbsaG
6aSqER/6nBaiygB82Oi4WwK+kRe/PukROyhkZBEDuWI3DBk/T+E419Hint8YL8pFg7K1UttLA97S
JoIgVl913dNwHwtvrPrF4q3mQKyOJWw/y1rCwvqWyTDsLqw3kk9cxxnQXko4IAkl2q43ea7rYRO2
fcBQ0fz2DnFuUa/ld8q2Bs+3d6p4P6SDn+JvxkDq9PyIODA8cZYpWLoiQa4cDTqYRA4mHD0QqhKG
KhhzvI9cNiq/J+fGQrWffRsj4Pm1+mztUAMOaC/jWLDaTWOD6sJsEbUEeLbPgPP5P8JPalWR22Yc
X6vi9H6UQx5/anPguRYceL3Nfy7vvnca0D+G3cJaQERTcATB3iM8GULa9PUUMvm7wudR6QK5zDbM
6RKiLLkzmdcWZLXyO6qcWpftSNHaeW5GQMYS0e8UEHrHO9oAsoyBEtmYIhjBdE4P5W55MGfMgBBc
UYIlpSJoa8wY5AZX8u35a/JNdlpzTQRR7s8QYlO35X7OrYQ1+D6Dmlrri6i79pPZg9B9uvTHMNYN
iA3gxV7l3aj4Pji6f05M7aXReX3nRPGaxkXe9HCS09K5ffERitq3lKdPtJ9fVfVYgH1ANMEgJvT5
J9r3dssIFekmIegPX572pmJKNaZC616D6zo+Iz2kFBUlMh0VGxgYY62tlmMEEqO5fdNOanMB8f23
VMEsQ32hyqxK4c1i+3UhjJy7hNcyio5J0+YH7RUzL8h3CJy3u7xc2icO4vWNK2kOAVCwY/2prEE/
bvolRnlUuFpOf9KfdPhrvkEF6L8daWwtjJz/Bd4inSq7HbxBBm2NFmTitsfcjOaldij1GqpkLTm3
JpoUr3bvSiBHc47hLA99WKLypKDeTqYSB80hgtep6rfCgWEZLu+JZIsJTN4vy+xrgOqbA/uAab1f
BtKwbMRcfhqHfNM6ZR0slDNgpTFre1qFVxqDRW5XX9JvcGIYzQekhXSxyJKHMV74nQiuMGyMQpbr
aGaHmbQjMqT/naBlng3kARZQdI9gg3z+qTO2Xg+WymBsSq/zG4tV3J1GuVyaetqwu2NUzXsYywWe
sK19/UIIWYbrjbc18Rsq3ZTvpSosdQIPdZhtvd72Io8duJd5fV5U2haWwiIBZwS8pAyI2wbYQfNX
CDbEYqRuKsUKwNraWu+9bUUnMJs/cxQLa25KuYsOgW+/t8WUJ7MY9f7sngIwptz51DBojDb7a5eM
J15+zllagB4SDoQbFa+YvYWeR+thC69OgvzFNQxwyBCrZURTh57nUjMvxj/q43mFhZ+jUDawUuqP
754bngB4UQY1pjEbdQvc6wpfBNTQkpTvcYoGvOkvRcCqjBkfvWD9YM9IvqzpzlWgXqvBCdAL2Syp
0f0Ct5fMQVD0I2VHi6fJCszku8D9YraOYRxsybUxl9qWfIgdYlesp5Refowlh8jGnGgJCYGQo1hx
yO3n8DOFKmMKNpxuDPjpyvq2Y97EtM1+wk3DkcISWEE1GN9N8bxMgtseg2tcWdKDnxR1sVMnUCRe
bFhTfZXdMhXrgsVbMmql/qUf+0yRFrULJsZBPo5RoNolPfZo5JfOM9jYVkUFRaS8apLfnyzCZadj
VgKWpS2q66QQhCGfyusp3GrlnowGpOe3U5CDE34KIaxiKI+O5jycPa+fq93NxCDEu7yNCZrBwPx+
FjgFDAo7Fqplng8T7c5Z/coNNfid8SFXiaI52jRR1FfoB17UPoWKasVhmG9I+PtH/VxYw++15eGu
/zGbgK+ySi5DhDYe97/ThM9pgATcky1ecinA6UgrCGMcQ3sUQeG8KisSI0VDZ1VMFvtdfprC5c6e
ReAeQp5aVhGOGaaXzISoP8nTTAlG2/tS0xY7anuRVoCd0QUeVlcdLVwGj2K/Ney32xDg9yno+t6B
UwisuV7YO0Gk1oymhBnH55dbJKL2Dsyljpt/7mTJOoYuU06yM8mgoTI09YKB9zOHrwLy/IvzZDTl
z848gxyYeCA+iaUat8NaZ5UCFM6Qcon0PSEiEUH8CVzpxT9+mOFoUb2Gwb1A2ya3JXF6xXw8/+8s
KndQwXuHsl2KatKvx4NzNMhdoXlrNHPJkU4nYxaMNa8VERPqKciQ4VaKBu6cy80xpy0S7n2fNfQr
nZmFdPJ4mt44metnE58h1dhbSu/UIldkzQO7YMPJrnRtjn5tW6aKlJsEE4AnIwFCqoiQwYy20NiL
+RVKPjVtIzQugcZ60em4Z+RIbg4U0/FlZ6+bO1F0Pc4yHCyMIVNzHsjZQOY1SLhAlkrZyh17Mjbd
Dsc79coO+x7nYJDwPaT0TqCfA1wnmobkQQ3GN3MR6uRoI5fc180zsZrxz/4AO867qToBCmAMo7jb
k+p5jlzD8Io/AxCHLR3QB7YrvGHMHD9vcVKU9kTO6bkbJwm2mdMsrYPHxdiodrxUrNVUdSPrjBh7
2aMPr//vSIcvWITc9trCOfFv5O0jLe0DUJnG1LoFGhrHuty9OOtcwFCiMUkSFRZucAfpFPo8yD6y
iGEZOjOIy49YMOc9tmAg4emg4VDFDzGe8OkwBNz6ctV1jeD49VY+Mtpd36HEa7y5igUkFTHugIke
wvV4ujbGzxYBKdIYQm/8RUzLw48p3rvUno4pJ/MCkn7b1++8E+P20tRaQp5gJRu7Xxwl2mLJwLTb
GrktmqmoY9QiaExhxnkSisJ5BL+niMAF/hbEe/vg9OFqxKfI2FAtMYrWFoVzVSAQicVb/Q1xIVtm
pFZZOa47wweNYEQp6jkdbUiUdEwlaJbHk6e9hsf5J6eJa3BdF6WgCXZlEUSQ9ZuySC9jCoRqIXC5
Y6FteuxyY2Z6O/H0cGfF4YsQFfjOLGCRyDpSTAAQ4HbnCU2S2puMOUypDo+q7LvA0M5jfwD8C7ne
6X/CMaAKrUuBY6JtfvdjYeuk9aDLIOZc8GUgjzvZHgGHZfN5U6VNHvA5s/hajCWO7ciuIezM1sLU
8gcvkxY9+LGW9ocU9qL0NJNY6HOegNOJL88nSDnSopWnRDHjZ9AwWqPewJpRoKbgdfjwG2jrDaOi
ARbQBCTn8tnJEKMEx6S6H8ogjRN9DD6OA8vkRVg/fLUBU0hrfXK00WhNb0VJkfGItidcQIY73KP9
gmK3QwXop8SgrMrjEohgL9qhLu4rrHB2L4yeoPAEfm0Kc0P2dr9JB1+eDs59TMhaHmzGQXeYGIeY
Pogm/pspLGXAszZ/f2nw2INOTMF9MGw5HFhDn8BJtJKJh2OpkE8/s4KqvyVy7iDqANZF9yre450Z
Ktob46zDN4bMlDNHz8ryj9G8bGIoxEJsS7N+hO90T9HRmdFQ5AhCO7QQcuuQfzngIhn9p/KOosme
y+SBh5O+zV2V59fJQGjYEjZYiFhRDQkbVzOusTxCsgRuMZ+FFnNfrD08RTfiTm2ZEzq14QZUhnJg
3WqLKix+hPXgnXNIPJoGMYIHGoOdyjzxIDh6xigpNalU2du8VASYJT2TM3XtG21VDYNF+AIoOgFw
DHvcSJa49cjX0PVkE7SHBa8UVCwc+/e1YjdEge9yH9WG2LqkGAecFc1EyKtPlVZXWXSyNIn1NIbJ
XO7EfaRe7Hixjr8efYDuzz6yDMaIOTUqcctG4s5UpVIoPyzw33VbWV3eiAz//1TTIhF2VY+fTzCC
PTQJKXpwdCjT2pNrek+KqQt3jlXuAfChYxkHOqhEVs3DcHHg8jdExYU1Hp5zt5SizO3FjVfIVIUW
Cqxz5XE3SPuRKs9fSOSeQQv9+8xTywyLY1Gk3OkwvFw68F19/qt0hYCzR1N1UF5bYKRw3r1b2cEE
flEmnevXtWuDFtj6T7FExjiKG8hLg2iR+eM3b9Zjp87gwTdmDVfxCrGeYtifOo3tOXsF+ekmtEqH
Zay34HPLqwLnTQI6AGtys6Hf6SpToFRpVMOnD0RH9bxM5T2Jt/aSyDrhm6NbU4+V0zUx4KsnZbrS
RFqkzzcFaAQG998kfPX0HTbAqYyGBBxmHvZcrrBOD6hrxPGJzazOPTaSn3VbfKXhQFiy6HBvcQD1
QYRdptlbyINV53q/lUrhvk0StvlqQX6AOjsSmFopSA01Wo1vqyQGTal8itSlN+cQNmEFiybQehmT
A75fZOf1sNaSG3FpzhtdMt0qcKyL7WJQW80oxO9a2TMwVbEIfMjecLM5pq0isf/WPd6czws1k9rH
Qypd8N91ruq1emq323i55nwB2TbfqKe5y2lNNVGUSFyaECm2tcSI6EkLRyo1aP6na+GESTzvZ5Se
pG430DVMCMzqEhJsRr+qe8W8/VWIyedTASyxuWfphHmwOlzb9qLmHRaSTS+xiNSMSNHI65txl4IE
wyAkpmOEAChlQmutzllkSzEvLPSZOhFCIklVkSb3PZvJTL86dp4uuQraPYh9pB/ctxvrOuujB15b
URCX8rY3u8iQMaS2a+v4X1dttsDRwxLNzIWcDOrtg6r/7bGP0xf/UJVTUoyarCxs6EK/icIetMHP
A6+MngAJMKsbeQYnTeWPjXtH95U8kYAYa8XdGO67KzmBGfaAR9hQGAh4b12FzWZ98pWwSDNSaDyV
y3qSlprEdzWrsmb5QybuO2DcaRXfWPBJNHFYLrn7HeRIwSywdet2TuG/BxfAUpBfYVDn9kFI61Ix
IhLGsjoJJsumTzp+xPBAehNuvBgf0eGNzjbgutP4+P/mv2VbapJe1fylEHfvqqAZtdO0q1P1SZqs
8+hoSqdoVPBChux2nPa9+IAJBxTF3h3o6mEettH47jDGuUax2XCVdLR2oENWPz2bj5+ZB/fz/3C6
Y/nZ52SEWtBfSS/Dn9fTnZXwtKuQ6WBASdW9oBzP+hHEn7//B04JJwdAmaibUovtuYXM/MiLcijj
Bok8II20hz1cv3uJqWDOJjgTg2KmaDHA0F9ZUli2wTheCBmhkhAfn9Tk9NwWhZNjqQgMNRYFFlaE
YlkZgO/fOuQBB2T+EgzhgdNarJD2TIImw6v/TfW4EbnwNxXkFknhecNVtl1K5M9CzqCv57TicgwL
p3S4cJyvHUtxkBhZTyhsgSL0rz0oWesrJg06P/dbMX/OU+24EpU0lqEcYfLut6O7InQoULazLWBn
ZppTkhkz+MicvSmuxvCs/wOuyt4bDUzTNT99R/AD4YXerOD1g0rYvZ7MC0NnaypewBg5FMLneoAp
KbQg5xOt526E1go0OlXK6dHyLwVh2yzBh3/d8o81iFjqdXrcZutps7Bqt/uElAKuDT0pdryNUmCB
i6KK07bn/6HAzi9o65bj+mJknL2gr1ZsPM56/C4Yue/F5OJiMGwWnHmrYK7W9jeXw647vER6o5Ee
rCHWT6pR3WGfLAoR0AtIFQLkEP5EZ0DYgpkgIQ8x032HgeARpiRp8bbL07oP3ycGNsnVg9MnJX9k
cD/xFobQH+/00EJ7pQAvbYrlN/mXHedpa7GFWoxO/74bzsP/1gdAWoKX0mFokCRj2WM2YRP6QKGb
GLQ+/+0KIwL2+/PJMq6LDptSqldtSS4uyqM+iGOs/xZPdOP6ANRBb3losMImQG97nPwoan1y7JuI
+6wPelCjRDXHUyrSiFUsBZJp9gvAYAWvMYohlm3ckELLUCXrc7k2mSFbL9FaBNwD38uNOolvcF8b
Qqz62LH7oaLHaOrb4vW0X9Oo3WKv6bSPiVlEpwNF2vaseXJhrYpRXGEowcaepx8pcGAYYmPrEhcN
r3etMKhy2IcdJYztgFigCz1hu//FHU3jYncld0ClJkMsz1by5RfhcO4Af7uZRB9KqfayAChQSmPZ
6wqf4WPPH/oM/wPr/atk/SGJC/4rybfRSncBEEWnuChWUTeY0j2lHhCfPdJo1PMeXtfd1f4EWBsm
f+jOe2I1uqwfKunLn2M5q/hNGcE4CL7hhUsTUMAN0dQN33R02ZxLEKCsCmzAkBw/UZdW80NIFSg7
1qRaJDoiUSRQyW62eb+4fdeLi6c6riCBikTogT91YlyfLaoRtzwas8S8bBTjgkmOyDz4RpgxSnb3
cyqvsF1OFCaITBUJBywAOFCEIR/AKPe9nHKbrUYG0ISBcnyb0sXijv8HRwEOW5Oir1ZJbusBB0HQ
NfDR3UcJmlqaLhA+5McGPC5ooE0PxjfHrkXxTRAgRER7g2ZtvwRpOlIVFvbK4UpS+HIFoJRCgzpw
S52L5o2uV6utkatbu+gxVYp5FQ5YG+Y7CK+KTN3nhM5bZ3zEoP1p8gI9w4oZFQvmEHSdLBh12ikb
yfCu9c0M/79/SMIXvvsKu3Ken5+MCWJq4FnlFgBPbeUgaPIYRMo3o/3NhT4gLjz1Oi6tQBwkTSZ7
8n3q8kkjI6V+RL1/4aMCi4o4I0Yn8naoZGdkU1fbpNop07rp/c5q8+Mz5/CXTs8qvpTnrAuk62aR
dGzX7r1PW8dvKkEPnMIEbUtGRy+LG+72aPghPI9nZ/MTnLWVIlP42xyzx5S5s+hIL7BeKNo/LOqR
+hM9fH+HV1noHgSyDMr4GgvzVTVKlI2XnCyhIF8/SXq6kHmI3sauU3QYWIHDujYaYvFBKVyBqTJE
4ZNF96LRRVWmuU+qMRuTZGnTnam6vDvy299ow/wkwyXpTxt0OC9U+Uu/E3F4B3Gn6xU66h9fc/wu
Fageh5zqqHKRnCwHREkIQFm293kZezkY299jpH2914hdioSP3oDhIaXU2yOMvFRd3GpUcdf7oEes
scEMrkA1WAihhG1xSYTDr+HQBhVdFp+d14mMK+0rpybaQxBwhPkHSaaqHbrK/ELgbBkRsxtHgTv5
K/5u09D6gYxLlD7eUTS3iNzGPxqUXbgZRwD9+yJ7uyB7mcV/xCcNpURrVcloeKBdwSHZiELNPfUM
6EpxaeUSztHwz/4Yieow9V1fYwly12axhPgo/KQGMAOeq5tGJlkF2Us1O0PdFYjkSHv92GI2sCdg
w68/FffaTjt9981P0c4Uw3JbWgylznfDm0BF7vfAKwAmiQNP/w+Mu27ki+wL+GIPK9+C0DSCGNlr
/xTSmf1VCJ90Ja6Cd6H6oMczR7KeXgYAoXGl+PAzX42DC60kZgLNpkDIFR+8jpNx84LvHqmI0CkN
i/8JFkt0Xo7qozS3IZtuqSNiyD5rPJyu/HCyJUPqMDEv9YDqF+XZt7pQVtC1eKjEeoG8g7sZi0fW
Ww8U7+SXfFOfLudu1L+ZjOO4KI+3sYcHkoYTINwMCQ1cgVqBf2FTbAStnEBLNJHpozt1QI3IOvwe
ceQfUqtYl/Sr2CZrO/Q359L+WTnEVq5tqVh1GoNcWLqm6z2h2UfRDPKLkcPL5bQgwpnzNYpRD9su
8WsYi0vMTZrNv+th2gjJX7JfXANIctwc/lY9rz1Y8Xumk20C1k1wn+VxWcz3V6OmgILeBk5c2QJr
21n800/Nc/Ofb6PC7Wr5HH+CyVdEOYQewrwFgVdpifSSHm56JU9SGyOIBcJviFXvKzqF76YgEVbx
/q4RBwlEM0YH7jRbIEe2GduUAMIzR0+zD3EcfTPQLIoDlko5ohxCa+y26JbSJd9o4EzctNb9LaK6
weWwPiGTlA7z4vtnhcZT14sE0XLzClPskHJuOdof8xkwZWqYTkjOcRI2G2VDMJ4x4Vd5vHQkubp/
6fHSbSgrj6qHEROVBMdUw/5CaZPtEekcm9gahMj13eEnifMmQe2SVrkyJWYQqYNCrpojg3V7tboM
azFFiH6z2fI2UP8q1JtXD3EJC9hhJSUgraW1ZqX9F7nE8VVjdm/b445rzJzpAbXvbMJrTgtKqJHw
uv2SIvx7rZ7PvAbhSa3EXvvKmRlOwvsa5MmO7J8NOOHu9yulG0qSgRs4rDOyZM86noQ1HWjrfUTm
BPeu+L1ELpdU4JvD6QJ6ArWqjmYeAvcHPgDi4ao67nmlNGR6u1+MtNUicsjbSCc1LyNBnMUJML17
7aNgPkWMyq7q+yuDZqMqdjDz0z+tFuE3m9A25LhOefh8Ak7MBOGoX7vcPlKayxjXUoykXzMKq+Id
s05YTv4CqXWFwJ4FDT3nhG3/8jyZU10ShH6t/af8GY/IzWuRKNDsHJ5rt6r3cPkaTRPPEwW8wFZV
5sksMACT4e/IGflqn1DNNj3adhB0EGMddc7A1Ka8imIEQp+MLoAr+17L6kRiVwbGAKkXlyx4zwXl
4CtTSyPgoYyykuW1y2BIf6KgBS1RWlNEGhJxmiPaCVMxzeJwl0ytk48ej2sLlwc3LY5OGiY8agVp
4rkLBhhDt1CCy6czTSr1anWC1QZsQ34tWBIekuJj0lfbXwFkBVnlKG6sX+kHI5H+9tpo2eMs8Mkw
qhqqbAv2t+BDWhgPBUBteAcemkOS61sK8PKZZ5opX7c8/2xd7h8Ws8MmwXZafB6oJEPT2kbLPpEa
aSG8TwJshFnm1hMVMLzrdJSTiyLhlBltEO4bC2eGBa120Vsd6CZPcqss4QX/JaxurwNEvQeuE5XJ
Tq6eH9yWENRyoKPh8AGfInnwn7qMZIEz52vQtlScNIpIIdG9JwLg6EdN1kHRLCniv78qQZjF20jV
fEub2mq26HANQ98GH9lyriyWQ2gTBNEprzGDhvK3TOo9wCUD29hndbHeiZWZYkfi6VRgQrLc50ul
jxiMzcYEk3iWRQhvTcf7vuEmGtpSiB3H+3RcW4LbjXQGl3ue3iKz5tBb+gLVUdgs1BVpkmrcQ7Ee
2sDI6sa+uhKHf0P0vB8va2x7OtGxEEqAP8p3F9d/vvc8eSvL45RxS/9V/DTMfAO+L2c5x+nfnEBm
BhzcZC0hJa81Z039eorqWQlcRx9PIVrWBzAW+Jlcw5uA2ZzWC5uU5YTSosRkAwYOUDGVPEdM8XZB
QcDblzCEmjcN4D8qOQfDwkOU8q27lkifCQ5AIU7alovWxEgZQ+HP+15A7s2J/dmnatTCBU9qlBqa
kY++a/iRUlW6IP4vqxZ9kMIltL5l2W/UutwxCKHnxAqykzaMOWRDuTdZQMJ6Dzib/6Srg4ZJKYMk
ib5JEs2xsbWtqX4Nr2iToXLPFUErfhaDDQUkDF1+MNsSmtdXRkkHjreqx92KYDBcirRIxqK4qZfo
Nsbgl6sSR+0ddbv+uHuE1JqwFpDqyqWalGBc8dOcw6oea98nkzfXJ/xK+q5DExoHBYHcS64hQAnp
jRGYS9hKIWpZAZgMk6v6ReVKqR0kbKZRBS01xtKCw06D5HBpgPK1N8jWDDk2mBO0vM8W6o459wUr
IBmy/PSnffUBADNglAKNx3fcxFnaV0DgLPsiHtsHbwt2DJPyc4hHjQ2VPA4XtgaZPh1aVfGK8x3w
ueUvANmCnkV+JjjehC6zrDJZSey73O7b/bSTY3qJMBcdN7ZmuDLH5tIwUcM7eX13ZuNXy2Byb9MX
am8Tddor2v/fDj2hpK7HA5Xt2HnLKQnh+/NiqNUCzNnapYujWc7HdZP8Ur67G55c5jzas9tn1rAw
jGO9P2eWZ1Sl+UuEACTsu0juKdE5xMiK0vXABgQ5HEsyTqgBBJCuytmle7UXlB+vPUQurDQWJ2Ro
uct5aBHgcbHtE1GV9VJjWYuDhij5dBTN9IOal3S5yVFZay5yVwSRED0YB9Thacnk2XSJe/buHXme
B2UuTHZI96l4LGoLwjGBiTA7KTSZFO6w7u0mggmeKPswsvB6PMIjJ59KVOUv/sQ2XD3U29NxBz4W
Eg12/WknK0Zr6yljQPnn14/VO1z5X77VqsEx1u8Gz5syqi7Z+3bRJQ+GAkEpDFemcj+Hwrb0GGqZ
8/fMA3ecP9M6DJhX4RnmHM+RdUu0vr5U/hYvMXUZ41XEKTG4Ang2aQfA1iVPwWFhKXfEjckxi3TB
6gIT8zuxKPUBXNl8TBBivK5V1sBuMWylyKYVBu1p80MMtS9/g1YFtGlIgejoWv1IdZhEQml/7jnF
UAXXoAAm3PDa1SmtFJoZUMrAIwpSnsTYNm+MQ6AchrHskbOyAjRM+FKPX3ONo5voQtOWHyUgF6I7
y8awo7Sj5Kz6PJoYcbggnEUElk3X+p2FQNRamQs1KzVxEGLZOiCI3rhwMktN9bqldoAd9mX+ZIXQ
Jqr8ci3HvHXa0hoWPlTuP4p3p08NJki1ETdQJnE53BXyDc6vVBoaj6bk/GfymsMWsbjapgZPGqDA
S22Cbv/DGMP2bXaqe7UX39UCWx8XkAuOs6TXY/f7hfFoSkN+PXjxzmNr0xL0Pdy87k0urJtPEh6Y
mz8Ic3MpbFnJde35MgBAp8evL1AhByDnKilHYC7kNU83XeeXBnDSE+WAlitfh7+1jbb9HUpC8Sdg
mWPC4MzG/MglZShU+wU190GXE/wApwSgTtA628KQ+IHLU0XPhCZfsSSBs10831Febl8FVkz6aBs4
CY7rBXaj6AT/EJp9VCnnyNgN9IQuFlTbbUzIdEYvIQNfwzZZmE0P7UThAm0ChW5/xueXbaF9FO58
2VyYr3FU7w0s/ISTMxP5zuqpI21SpdvFtgqpP1Jid060DJRaYGSCNYYkCC4O86C7EqXE57ExIuu5
132/58j0VrsP4rq9hCKcH7Hdl/ykTjpPz9hxYSd4M1tIhPBXwJmO3cf4JXmSwLGzGByCHjf2Ntk2
fC+Pwj2SxSN+3N5yv3i8LAJFLDFvPQDtQuGeLK8lqR/OsSYvBJhbgIDc1NdwJC57pv/dcCOC/Z4h
SxqR3Ig27sxUzRr6dIKg7MZmVGlHaNsS1u2LtvXRbaii6iwDGr2CyY3UkZfuc6GH9YPOg5S41Aln
iMg+iw8uDdXjfLcUaGssExVOXJQQbGa4V9IiK46234f4REBpM+47egy0sZbnKPgIT0JIMabXu70o
8+Cp07nBk5+X4aLfRrJ6+DvZr+GhZ765aBTw+KDNiI7Bcr7pGRGZdIs5m5lbX0tR6XUBSEJIMKdz
VMnfTcuDJtClSfNdwy7qNUUiQ0TIKc3NU0VTu6aQPt3SF5x4F3geNAlBIsLhe1qs07ScY3WN1iGo
PdeUUTxHiI94H1HcMgd+8cOlPDCUjstqRn/ItgGHBIY2Xla5mTAn2q0R6V3PzvmQOkMVxCJLT2Ar
zdn/bSJsLc2i1x5YkR876Wc7rZ/BpuJ2TbmQbwzCN1vwQcuTBbCQd0Y0/w/hfrzPdedZUvX05byd
kAGoCyjx8KOeUk540pFOCzqwK4P5fUz5TcEozsSFhBrmtLZRIuh36R3bJMnzFLizvE3a/R2/KgoS
Sll+9Jo9GZmUUpr2k7JnzY/Xcslw00H61c/4wew5oshzrKEWp1WYZkGzisJ3mxbERL3UpGPSJSG/
GKLF9xrM5tE5ws939XkyAW0BgS5xmR7X0bjqhouxyZzzkXj5/91e4p4KE+E4PIGx69Z3fnNlolIq
qKV5BkjAjbLkWOVOypkb7jput9hXcz6qR2KtV03kxiaKqTwPPDaxiivMWe1fpYpTDlhWsw8A455q
aIPmh9cuUjolQkQAe5Mv8tiko4igIkddZbQ3/71OLtwIp6ZpXsMdv5cElELUzRGeZWiTglqmNyWN
wESTE3ig+QQU26Hbp7euKPHN9QwOQI3f+/KCXcTIekoceKzp72LAhG2kK30xiuYXjqoz6xYjpbiI
W7eVn9GxDYvVCZKXXRbG7tM7AoWSTQYzOVrHaTwy+6Af7AZjRpJVSNq0tHX/ljVuXHTDwb6vLXd7
1yzJM2QUY+S7WFV+ZDC4NKwMrO45FllknPcSj8Ne5Olrzs3fnAZKO4SSpsg4buNoqoutqDSL43Y0
TQu8O9MbCRMCRF2f8HNsy4ZOGa6US8GkB1qDDB8B5lREdYSqE7+kPoRdxSCzleh3T5JrpmWVBLcK
sut7WyAD/f7f5F5nQy04aCI4vKmzlodpBDHJp+UkmV3VWk65D4xTkV8bkiYwZTFE6MH03fKXbdiz
2uWfJIBhiJer3R3MXZNBycz4eVScEdKVi72m7mAbBm98vN00znA+lsxKWF/dHlTalXKIyN3VssYb
oORItf2Iog9JMNxcr9VDsD3nA2Gr1vG6LFkQZ7NkB4y4CstJ5sn5syZIS+xCtT2iVYprys+SlwT6
bS0D/qej8teB9wfO0Ivyq6YckrrGZTkduxObo/tkT/aRo/MacTtil5YL5uI79aY45ONEZHc2G00P
oq0Oh3815dFmvWLAZQSMeKJmNDecegFVsw0Tb+CGog80uQW3fBPWD40yepj/MC/15v0fQv905dmT
wDRHiPx74aaVG+QXBsiIG53pv3ccAy4vLje+TZtaDPEPXLpITnXpubYs+x5ZXGI2oJIeMn+6fwUe
T8SoCJyP8oXMDqOSRFtAmfD40BJyWOQTAwprKEiTuHtbvF514XsRZY+shiBvfEUFqflzOU0BmniD
vduEy9hvedBiS9fYNm21onrGlwdNR/lbNHk2Ya2JjOqXymY+005eaXTveRPPcQ0LwEMCo4wAaq7W
FPI6NwiUfxA0IT9AAmeFR3G2CsLuqLUDnT6XCuJl1k0AHvDbq9LlNsjohE5mrJPDgb9LG1hTdSlx
ShEPR1BzLJHl/qAdY6In9h5C4dHpLSIIhVgEtGbiaWWgb40StZQk3vrjPu+rHAq1eCROKZKZnQSO
0hWpo1ojP5SRkU+nvT7iQ6bhZxcCVRDMVvjgfN5DYeEBOIO/FzqqG8CIu7rNmsxjLxnNlBI+CnTo
Ywf0nFAPQUo9uUJMJGLb58xNcqMRbCZH7pIPDRrZJeksuukqU7lsyafpCi0I7QKTqT3dYRM9vJd1
PDIIDdZdO+hDP3S2/Cu8cwOWryG3P9TX+UjtslG8V8EMVR6G+blw0vuUn9eUZYL8pkJsdVO2Gddl
CwfBI+a9kFej/ZIj/MLYk2+Moiks8VLaSE5hS4hRPFzvomDBPHIuS61eiw9tABrQwDJqAk9plKS0
/aXKYtw+z+/05lm8nHE/WiVPrzhTn7KkoTzGIIa+IBBLgUQ9naOaLprzUgTi3ObXxmT7y9OXKcdy
dAK9xVpO2WUBZQ0lS/hgbTxJRRffmgvpv8+ADiMqTUihwNtXrmP/djPgYXJYt1Wn8E7/5cs/sWQn
sa4TlmSeAuGaf5AgGP1420FOkb+9cLNRdpsY1/puztoFTkJ0HJBdRoKNke3Lx5CgpZ/yGeDflXmE
M+iGb+tZYQsU0/fpADFp/qO5mjd9Q/djHnlYwk6RMyDzKAWsV/Vp4SeWzjZD7eKPwuHRY2m/eRfP
K6qXbGU0neA7YqDE8FAuanvHUyMB3roWnp6byEtspeVre8LnB3mn+7M08VisCV7vNuSuq/c9K1OS
klQMluJjPetJ45zdQU/+zgly90Fk0EYY4YPIeEQbujfjDM1t6egq0IIC2Xgcu32bv5IW/OakrpH6
YwugeszKv/fRUvrzWMTy8pxfcHspXMr0qUTFNZSZg2Sxt7r1GLL1fU4p0K+LHkolB2a0BU6F7g4Y
pCwfnlcdOTF5KMOZsUJp6JYoU/c2L3SJsP/OxjC8M+yPZRCWP/D6Wpp2EkCoRK6AgMva6zuqeEDT
k/KMlvUML9I+ihJ5ebNhoKp1hZwCv3dE5Nf6C2No4GnHBEAVWI1DPrQrx22T9ZkP7ZmYfzzizAff
PWfHhRz1kneQHtr7uzBzwuiojmjViLFiC1rhrN0SxFMlODIQY5QfwmxMxSj0joQnUVqM27bG4osO
atg3m1bt+3Jcs/ZP7+VgA6lULcOaFHkoCE9Bi6RPINJdTsO2MgFidlsSMOPqrhxsatSrrU/yv+ot
ldccH6I5BcK6OK3FXGhUf2YpMVNQy0ldc8shBID5DH2r5djjrApNobbZGlUIMWClA1oRzcacy6JS
wum3payhg84ybAKaL78ZM59V8lOUmdg1a9xMHdaaBzp/qkib6gu1jPhrk7kgyAeBSuEwLq9WKos1
bpxYX6xLKkb0JggMiJ++/EOco3iyUR5GFI0GyyEhjuiNuBjefujxtHTKYi/nCBXALxA23sAheUHh
Y+fQHMBfpCEUmFfEfxt4YEAXMqPhldoB7CGri/S0PPVLRpCIhyU5z+/2hjgiTlzRr5bbRgXOGipl
i53/3RGOlbv+mnvHmPynSsjU3susWX9CsHT79HMRYNKUb0zeCRoS4M0VpwIkqNITIaEb2/uu7sTy
fAElOhruuME4JnqWRVtagfUY7XC+kmZjjU4bZKDJXb0oEjMEOVPPSRlshU2d9lq7om5hU0nce24l
TpbJfC51fW2MFdF0d2Wb8tYeKhL6xgf3kSurkP2tUryac/6y5rs5j8zmldTTmM2FJcum3VqkyKHW
sXJ9165gjRP2hCGkkqkxkgLlsvfw0YHuvWm5ocKg00kYnPIW5RW88zt47iJ9hKEix7ROt5u/170m
zfvcBJVIi+viPxFdgwgMQdb+PbEhDlnsM4N3NWsoFPPN3DoOD1whSrRhPpEr6KyeaPxHSLT+D6HH
3WH500QECBYU3Nbvy0tS5n2E4OXhHq6l4RSwhUFvzmPEONoGbfoN1Ca+7EKDtt6KNtQY1J3FdWSl
pDsK+Bq97u6fwqo1dOYsL9VvQWriNY9JwE8RLb/QtNxCy6RwXcu0iFoLknuT0AjDsTKrl6Wbqpsa
RUnaMBh2hnhG5ENlocdMEGgDGrVcIVjsL51mLu1cWOagUTJSG/LmnhxX1wF2j0pk/kq2Qp7O81P+
kqFk6CoM+1zUIU6BO2Rvap+ax2APVUCwvToNn0QeYea4Sr+kzw5/bcdctTmIMJip42DJuHWh6l3s
xDHla2Bj28Bu23ve77a6+bcrGy7Nim6Eo+l7djEHX4XoGcXIF1L9y9L7cixy+7h2qYm274kn4HKY
EmqYGeLtBAc99ao937dNf0mtNcnIcsba+YROCgSLRWOLnTaGoHRhwnA+sqtheM+YNmNBVjnhsvBY
VV3v3DJFC19fjBY5E8MJJjnINA43bqKT3ZMQRMOVkkg3SOrdm0F2jN1MtRRzHA0lZjitF17HPa2D
cgiXqhmTjZrKU/ac1p+tmi8gAMhBYTbM4UBDXuTZAwcAmtW9GAyuU06LdHdKqQhscHtXs3jnDip9
0RnNpECKi4NbngiUUJSilT3Kwq5KSNHJNSC5SSPMzM+mZk2veVCrF5sc7TuDa/pE+iFSnrEWtZ5z
nDViYVZE/XYaX2U/mTxyYq+hGKqeK2nCa/JY7Dw5VUMsX3ESVcZpH0XLB5fYQ/JHaQ6pTfHYwiF1
Ec7E9OSuN073mktZcof9PcWWILdPvoyL1l73h5dhR6cjCMIBJC/0FdwwNYssutPtNRELl1UvDHCM
hexX/3AP3xoy6HQzMLhvIsqRt4QSh52TWugJZiJRLCOWiCyRer1bcaLDeouoSUYN2uCL3aplRlkY
xEzRk0j19xJV+QvlEb5MvOiuZwxEjJbQXUHIMlMNx0aFcifTQ83TU4raH29nA9r0EHOpNuRZJ3WZ
f83kkb4KK6vpNnbw62RPgtkWpjU3UXzjtD8wmdOWNJ9QsHkxo35kn/EBXHPLZ5Kgr6lbEFXB8zn1
KnKOmUcTrL8UrpbWGg9dUboCAeFSEUowc5syG5N5e4ClFyC5esjDCriQ4F6zOkl3aeXQBgmsCBTv
TXqPyPSer6vuV/8h927sDNuuXDjID+vkpZqAePPonhI/jR01HtV4XTqajGdH505jSxzeoJkHtvOQ
bwfq3xicjATy4FXstaU3r9xUYApgBFZ5JLrnkZPqFbvt24jWMNXukcRQwf5JbKfHpHuz50ZgQ+FQ
r5jfotVINRoUHy3IJopOeslcgFgODL1bELfosuH8mSldcQkAcwvGpAMWQS5lt7kO13NKtwAHo7kE
+6vMQwz+2mK9j/bOARqxLGKWqTjuGO5ukz0Zi9MeRIf7FkE8kyeyYGLhEgY8gz/1yOxDWrOsBNl/
m3/pfixsAAhiJPUFwFfNRFlhmGq8BY+AZZXt7f6IcmB7rfT9Ac62SQn9uxZ3GdUJEUuysVJ+7uXd
YX4eQcdtR6fFc8pDiu+58mSPyAo2gpb6Zzd6W7hg9+Z0NYrSHZO749R/fTz6WTuOnYj8droMfy/f
lfzrq+OfaFm+gGKR27iOayZ3fQxr08t0rPS8lnSPxRTFdlTgVa4JoepHyyXHiDcvRC1UckLERnGx
PwSrF4VodeJM+pqIBuo+pgXxAE4GOrIed5eLZwe4UodyN47N/OSrEGR5AI0+pi++C0cPpedawZon
LF4vkT1auPsAdFREGv79CxWzlf2gJUI7/kNnkaqD9H+Z9FBHy0V0I3t8xKxzdCTinNPWx9A5r56g
8KYCwlDsfOjNEuAN/AVu3PaWdfiapzyl8RbxCjkSf9IMZauBLaYFGEXcNIJyPd3gQRcC0biq/uhP
HFoPDVDhD4cLVeT6gpKe0pFSsZ83/s82VhGHAs3ErkIFN8pRazP/Cb5jR24B9Wap2iBdK2GMwZzo
ET5JpO6ccFXgCMtY3+tnLchjEYwxzfJwr1t+Kvhf6VCCaXTnZwwprEgdk3q4Ip1YqlilC3axcFow
6LTo0qfeba8640iaX8r+FryIzuY6C20jA3IGzSo9ANEwjqJY9UDw1mF5ej9XggDzVlIJFDjdhEmR
jKVNtbQn8plVJmCLfej5qlZSo66awwws2+fF3/BVYA9nopSb4i+yEqKokyL+VHyMo2cIgVlmKVKl
P1SOfA8vAEyZ54HgZugieyWXrFuqe0o5be2HVQswkzT3wb5/e5jExeQApQZEy4yOT/2tnAR0/IE+
jwG0vagG4MqunbMPQWxPRlZO466hnEJgqrcqHylYKgTG+5BtbijZQjcJGT6fwwxCzrJ1quu2MOUO
2jT/FJAhB5x4uX5H5FdyawUfCS+x/uhqZZytM5EGh7UOhJjNO5stE/6SDStu56KDAMukSndyquzu
FbbeYvX9tN4rm238RWq++TutSnV8TVScXpy/oOlLlkpXdzhqIgubEiJZ9XkBrp4GO9bzNd0VHOS8
BylHKgJVK0BCaj/ADA2fnrtaaGmlq+tF9bByNXkEIZ/dbkfC1nA4oApwmU6dqo7oRziah3R79h7j
0SHc59px2Wm6sY2SlGh2iOzEv/5R33w66kkjlulWLPZCwJmUxEaF0SBWBVoB7Qh6L2bYrATyJKyH
747ROv9wuACtdc8xZE18J/Yq5QssHbzqKenyEVxhzIzlImB5vUZo+arWppMUz6YNKKLdlbyT4z5A
Rs+Xso1UKBk0TZj2deGkeISUaeG25/UfixEApjY1bo0LC+tBXljWG7ds8XFiq3ayNmUX8gczXx+w
jizlbWsanE4R3uklmGPaobexqknwqthb8TBN/viA/WqghKp8Rjj/HX6AV/GGpxGD1kdoRhfCSbB8
b/yGU0lk1MCn5CANDZb4AHIftdLAD0HqOG9Tz37LNXQMP2YH3EerFNPoZF0HHp3xblQF2u55Lf+e
CRLFlmH95b5DdjbqnM8Lz1vp6DCGrJ8R4IeGjHM6GQL8WNw3IIRbjOyHzdtR1hMVBlK5K4EB51JT
DI4q0Q3eQBcfq01oIQ4pQnKwTzrrvaz/qQrgA73DomTjyi9sIFo53vc3aAsASDPspd7cX6hGKNR1
4tHhOLsfM7tCE3SEDOp9h9BMnkYucmcNWvM84NfwcIE855R30hQd9qazV9O1Dh78+cG2aCThCuh4
ebnLfPbIyC35Er6X0jRdNMWjaBY+ItvHSQxbp7U3/G3G+HmeHTRXf+kImWEYZXxSc80+0Qg/fVHQ
X3Bema4DoTNq5AvBosNM7skfbMlbrc87kZkpN7HPOnPvmnIhGqgQFKgRk2tYB+ggvwjxnJTrHaVI
ougilO3gATpMI48S1Tw17pKUOB2W6A6p6MpzlLkFb+eoVFiFOKO0/uWkObcozW+eZcjzpTetba0e
q8ZGnN+/S366h29f6gB2Flm+g8rnDLFzGhZACt8eSIm++YBMWOaarjc/0uFTX606bCA+Iy2xDmQ+
TsdG0ykJWdJTSy64Ss5s6G/Tdxb/ECKQdzSnZwrMgbHYezqILd1V6q8MpQ56XPtUyBdayZgeN7xW
Ij5AhTGRdpTmd9WvjiKsAJFRxLa2X8THtlZWFNiMmJ9QyGSRHIxanF0ebioTbZESH9AGRXyxLk7a
sk9XKQe2/PyPhT8Fn5+3RIjmTcdOgJAIko+zTokAUlWxS2xdfCNGBQ8DPHLbLYJT9Kefenb/jR6y
uyHlyxGAQkcDOwhlTTTctiO5dBgWNxuz1HSK6kZj12eEfQIOfsQPBqYQCH8g/l8sMcm3GIM8MKfP
uN9J4mTMdhWFcVbpN4W39I6MTc+knvkgMF9OClbLwp7svBKt1ygWvhIcXRg1kpjuJK06OV20maTh
37UkDBb2M+O1OcGHmWsmsmI4u2e/81iNM6Xn/sQDq2wGs6VZ33rz2kY7MTaB+B4J1jgVpPfA04+K
lGbpfSOl4PeptNBm9Tg0+6P2FCZkWHX1gHVHumveLcgJrA3dr/fk/gz3+e2iXUWZkAS4o01McJdQ
v8c36uxxpj7c0Bwg8SFbX5fpvNisD9UIYLN5dMnISzwthdusSsT77pAJJKe9VxmHpEQ1h6j2LStF
SKc/281HYJ9Xc1KpuNwU1aEtEX/RWrdICBO3H9nkQU/ArVzBzfXM73SJ85ItpT010TrrQ+3gkX5z
BOJdPNmItshc+9oP1ilrhr8VfZh5h3wYQvdX5ErjNJq4el/zxJIUa6N0il0XgwIYxwTZMeYy/W9u
2EiwhHyOFulftFTxpYlu9Zzk8nPMpdsvyyTU5tcUp0NT7nBe6A47uf1cmqwwJw6BlOzCrzTi05M+
EqGw+9+UC9Q726jK6ty4eSOj8RygRLjWFt6OPtSuMkapKnM6nJ9dB+zqdGqZwUhrvBQW3AIwVs7T
OdHwWlYg5/KIeOcYbvRZHZMWKSqGJ7Hy4i/MatjOp0kQIhta6fdc9bi/Y8xGWsY6nzzG1MELeRPG
AXsuQzwUOvz/AqiKwnuP/aTSmT/0lHqTi4lQG8coePp668HY7qH50i0GgEoD1zlRYOAp9iEEAMl1
pacCiawBNTxJ2KXaEtLWeSVSCfSv1kVr8pQD6jGpLAmwrdaI4ZJNOi6WOqfO46l3cCa7etQ0/i55
18xjvmyaBCz2zXx7cjNi7hwvkftWtlKf/jWR7HUSFH3PtUjAStz0wCg+ot9b5sizbOBAqCK/fSuv
yMtzOQTWGpIDsGFwasXAQwb8JT5ge2anKtW1Dx5lxLGqrSw+V7GMMgUWmraM+BZdYYefK7mscFDL
8dUQhmUl1D8bMZd7hVhjABM1uf6xvdU8fPdpSERPL9rr4yC5r7ASEXUoE9IJ5qml2f792OX7rniS
Qyewsf2JRq9nYl95JIbrROMIe3nFSKO6BQHIPG4lR9Ywfh+13U4lCEhmLQ/6cLgBRF0+nqCeYQk4
8X0LiL22LMSe7sJ+/GNyWryilTsH32fCG94e1SAdCt9bjORpzq7+YI3sTykDS88wkPKczZDKNw4j
86lxiaAIwYKJSMkSc0HUQj44QKmqfMpoFEpolN9T6DWqQX3V77Z8EGGdWxslvPZ9OFswmuKkxkzr
ywmCeeFW0QaesJvIgyw5lIfc42ICfChb57X9SMc+0fI3qPgY64ID1mfY7Wfb9UxKLhkpzpfagYmO
s4O2YpydjdrgLK4eBL7AzmwAHF6erv72hMmH1mTWN1j3sKocuY01yyVnlU2VcjKesaqO8t6UGSPk
JijGWW+bP8Q6UES0fc4G2KRpWusG5EAGtMrwfueisLSlzcIC8gwn4Sq+Ja3ayDRhVv6jtCsgiPwd
ZNHnI7WuJ4QDp8iRvYiJazl9E/ZO54pnjgb+j1tF0c148UWgcZuQOswPV8Psy+kzuFZ0ietAZPtQ
WLcKMDhf47dk0MxWcMxvg2HV2Bcocj3XygSiYan2QKh6rwQi5ugZjktRU0lCOvB6eUnzRc/BAWju
ss5xlakgxxJQ++0THl/9CXD7fae5B5ne3lXurrJXT6h9KHD9elZUU/QuD5/C4HqICDiE0tp+KzNK
RJqnWNjXEv+kOiwYtDyUZ7O01Z475Djn3vVTlsGFo8BrSCx4MaDNXVfIZdKoW0RYpxWlt7yXh6Ls
y/xkz/6w0hyA2cX/KVOq3J45eY3kduSu7O9vgueNqReTQUCnneAIXrnMGZfsUbHEVYaT2RhuM9/6
cXsKJAvuK+rGI24s36pdaeabnr0yAQOESOfl7sk/ChAplYyAqlzLcnkdwRWTcFEv7u14HDaj4iNP
s+xXP7nvaOmxmjP39oGuICLHX1v6M3d/lTdIOF8qHbR2eDTxiGmtku0/GKFTdWxvmHT6I/1di+2L
02n5hZndl9IQrcFk1VAda5caGlQOx/cmOvdcQBy0FAmmzcsOLB57lbcOciPwWleyB9uyT2pU66nj
xc0lbRHv52qYslZZBjoPX6o/Xajo7glfcNxrp6KJx5sGaD8S4O8InCHwjZjeGwvJS5XQNVrheXds
WE0mGYD4CXtiqIZPLLMIu0XtA91PmhcGoDx4+L6oYnS3D4LPJ07tkBg9laPB4bmTDlmc5DBmJLg6
gsjWKPKvbqUUbJHFNn1EAp3JQjWAXFGaWhnh/UdMpXpRFDg4RpHATocwbTBkJ8apxNuJ0++mSOTK
ReUfoIs4uqlHYykZZYAuevZ5TraqA1q6h4ART28XDjT4kqBu5W8TFsSnbiSejdpKSAIbz4JFIZ5p
3Ynf7XpmxcpMXY14tZ99LhR87Vo22jrLLPpoXUAXtphdcYyNYsA/NJpDJ4AeuxNY9bTSdxVEo3Q/
en6IXMQqMpYdyMcokZdxgAifH1TNpe5ET2pe2VDdBGCaBXBi1BYXXcpoi9Y0YPTcRVfhgzk7fBr+
ejvnr3HBm6GjZFaKZnsZHHjDBhFiK5Ep9fqZKYANVyPooPq22bx1BMxrDZQpDipl6++ui0aGpmKZ
1EBE0GATrQdVMVPI+8pKT4Qci/i2Q/FJDNYC9iz1c91jNCZsi+7u/tA0bP5buiAvYJOU168kGC5h
ZkAEsni3rkOgfYFMsZiiJ85oAeiXRRK9kdRwSboo3yMLadLVNEO//dOHwjaMRR5u5uKvFfyxvMkQ
FHk5y+lr8ZSu5LpBEICWhhdnb6KU817XeGGLOjmN1DC/7ALx/VqFRGVTNC9XN/Fc9+D+i97I3Xp/
1VuMlp+8QweSLv5aYNQlKj0MgLboiczdkD6uaANwpqSBE7Vny30qg/VEQbkeHIQQxuWa1uMuBmdO
lvW3CIjPK37qJKimPZyxfVc7oIjb9FBOFesdHWcZ0NVSMoeh/mbvCCqtrmGBe0XhcANhfXR4YwRh
kK9nHvBrw1QQP+VPoojEHAeCs12z1szJopVEV75+9CzPTm7Rk4qs8S42K5DnKtybtyEraEikXSnX
QjBQ6aKx9zGKO/xf5zpoWAdAtCCyNqsSog8KGPWI3mD3AB4uLAHhTqtkCBIBMb9xwUkciwpVsgi4
oPo/bAgdeJRGaBp7XxduPUBBkzzsVhAcCIw+Aqrj95GF3Ap0lHTDWVX4LJUqq+gu0Bvn4uH0Cj2G
fG87WfevuQNIvKse2L5Qa7OR5he8wEUctMMUI1vAiKv1Axyrp40cMLyWSANtPAkCRBPC8DelcYik
EEnneXP4LvriuurhYAUoofxmxVQkkFxbKxe9dJ9x1lhCSkew7JjFe1ykOhSpomgJmPia/5/4HiBJ
RMsNBclQHUqtUJORb0zbFW1MpVRv71ThogFfmuSrjwkXUbkm1ApjS93OFrm8c/A6yJlw9W4ercvx
oMeWZJDD+u4mASCuv4IgI/9G2agCLWGguMWQqe9XHsT02Axsfu3dmN8cAq3uiAM6jxsTUfcXxunI
6B8JHhsK+ZzVTxblX7g91/H/cNCTp7QVLEwoSVC5r4/wQe805/9ai9KaUnOc+Bdht7HLPdku8h+7
GPTY99qEX5HQvpHQmA7qs3vPpNJRckjTmmg/5eOawVEl91il6B7ilY/wolj4QaaAU78ehurlomzl
YECgAshr9gythpvghz5aliREIrAQBxlaJ3prRo3IJadYKAQtl2WTQXJxklL0bZNDioURCp5enxs9
qdzOzxXtWTv/3nMmxCV1nNrk3rQx9WXJyzPhMB/sR/q6rKPCbz2Gl9c6r+4DYLb8PjsHfTSNAKDU
Pqe/I73aJ8e5tHuQdkqwdNvA19/zr8V85NlrwUBL763D/Hjgiu3kukRpqXVI56mEXvnwI2DUf4ju
0oqGYwT0mNVKuOfdAtKvraOEjRnMKb96NGvzbJ9GOBhBG/x9yzea6m5xPus1iSZiEi9cEHZ9CB4O
M7+1K6Ce3qjnir2dsVU0WvXpVjONkar8aiupIlrGVDWnPCbBJfHFNk38XDt80XKvWTgtjZU0YcfD
NaCXZmWWoZ8HL7NHu9E6/ZwCzvgKFAGXcvUnGBTKSCygqbkw3k0UFPlmZ2tlINBO+KEorNnSRcpL
D4dCaYAsXoeC3R5cZ7jl2536CntcVnCtBlUCletd0QVeI/y7/9nSEV23SRG1315fa8f1Y52A15hT
cPnML8f1CIyMASzZHmkj/vPRQOiG+Juhk36YB/fjx6xZoeMQKNTjW2EWCYseVAbQyOSsuNqb8vXG
uFGSLba7Kc/xevp+NtwVzENh+8wITvzQhjGGn66Kn/t60TuWl+HkAXdRxyczKO8ZrPwCFrAh6siD
d5YFwNfSlujA3QZtzZPS68k6lMA1dsKN4cHDe34mjD8MpEpSs3HAgY84FlTCRq6mvCzKeIkwdGC/
20AjDnB2kmx5IkjFM2nQBlDPg17DjOcZbL322Si9Ia5oqWY24oFuTvyPnnVnhlKbnmX2ktD4TWK3
Qc+mhU8xdv7aWaYLHEjJcD3GJmhD8dnByCniF0siCPaAXt2jv7DSX1x9y5gN0nTtSWGEOUdVUd0W
zN+lWIZCoYlUWWJ1Y3nrxLO4SZZ2uQwzbw/Xb09IGxH94QjTBsBBpKfyHr5RNWpfeU/y/K0d3KNb
lkvMYnNDMCB36CQLvFxKf74pBw8+E/d0Z1ifUYSkqyVXWXHUwodqD68V+/iI3+O6Oq+4u8LphOM1
Shbboyxi69HIWNCxyqhgT2NkBMdsJwx0mTGixA9cDtgls7jZBAoqspPW7yapF97cSCPo94b2fa+e
slJdSvirh9ns8aOjmhSXkozFmQSnRf5hEa42t+fYJZJNYr6Gqbk3FLmAtjaetBNP0YwVDNn7y3JR
g6FFwngX+cPHobh1TXghTPLogQeXfQJP6OKd4BA5KtZfuMrb5NvmE1pbX5QPvMIMqRkRneApua5T
Hz4dbVQbI2B+aAoa33kLlKYopSW4MkPGk9d8HREN13NQ1svcYeMspj9Rj1a47jqT3rt1e0YjZYdt
W5pg6Uqmqxy24njHpP5LrmhJHKPVJmgUiYtHFYRAEwyRwvBFSlaTkCkYUad2NDSxul6XhvwLmOfc
k9Ftd7TZubqJdPa/8YojIXhlfB2Q8Qwn14ZEUdzxJ/mNVyj3MRUsdGEBYMYwGoZ0T0Jw/ydm7OQP
J+g+tFBX7trNN/hhRe+DnleQxGEK+aHAfjI780KmO1KMcaF6gQPvBfT9yErRWAaXTIn7vLHBa4gV
4NkTOp7cUyeiRT8/sXQDX89zgQeSoL22TF4Qetc44qALuBIlPmUUVK921AzEE+9Ts/yrPdwNcwl0
4CyEd/lBHqjWteZLU28xxBD3e129d+OuQb8c/Lol7anx8nfXT9bYySGUoI+Buh3FAxuY+JrONH9w
SLc06z6QnL9I9HvmdKjqj73ebOSawIRuxrqETgEtOmPHAHBvCrIYRFkXc1omHT9alWykpv0dHKPZ
OmbrXl3PL7dgLI51FBzAId9s8TsknT6NB0a/n8KWmNw1kTHQChjeShgiJdb2hvH4IJV9UWeVfwOg
7D28O7egHvOztbhY9LRRGqjSWmvdsAgbLOfDyO1SL6TWu+ysvmSGB3rYlNuwVXahjLz7EgKeZlBS
2cmyk5ay/uo2ZHM8HpWkA/0RSoy5ZRU4iY8vh6VteJGpRTPR0VSSGrPlHDIP/2LoFcPZP3wWOr56
oXA33iXgxIqJnncqA3FiCPD+kbpfMGCFUvMM8+hJ6V8fPGYam9yjKk4ZUHDHvaRissQA6gmsxkgP
6lbSls/0NEtptbnFDLw88U2+jYOo4xgygUHwDiqorxEtimc60pEQtoPmTjYzZjx3UoER1tUg0DFq
UH14ybGeIj8qYPEubllS/5Jdgsg5s9Um1qtcyntMwZu789ic2juhCXO/ZKmhFbZR4njaYl03K7kU
7HlwiRBSOwKWpAxIYhRoY/GTsskmKkC2xVDgUY6+xlMnE83o57XG5bcLyqPL+CBxwu9zWfCKhKQT
DKgTC34+Xpak5yilJw6e18eJPkkhd2mitezj3uM3JcAB5tVH45JJ20+AruIx6pRVEz1r8Ig0lfvq
ZUfo97UOzyZKIcz/wcW4USDo2pPZS8XTsSZt2sHT8Cd/HsoNH5kL0xL54JMAIBq33wc/s3FBUmm8
KKZpR9V2v15NrEib7Eqh7aV1lAYEXnA5SOWDpeCxOb6u69e4sewJUhpmWhJTGueXDYaodnzt+FMK
Dqy3HT81oCUP+EyDbD0r6n6hnwF0GbzG0bS+gboKRDADEIK41R3dAnPakGIu/k3vSHARByOhw9v8
xoehgCa0S0wVSGraSsJXp416cuDCY0VX/eFC/Us1xV4MipNfSYTenDfldm6S85L7v73kkMHsjzSY
W1+Rw3mGKC6/5h/KAOv+J10r++DBflUg7glORG8gdnuwEkB+jMqNZaB0CFtnR5wNKH+5gbgsEVkS
brHIFVMOCA7GdE90ljzKyWDCe7xxkMCTWLvhky9o4/jMptwt8wMjPGvsVLmYAji/xYqKcOmxA0Fo
Q4xAE9S0T2cSh1jBA/tJn47foMGTr0mWYfcfASH8Y4chMi49Vqp8ENaMNjlT7CQrj7gbF3nIKOPN
7/HJsP5VywE/Ulb3BaoSAw1cMnmI/4fZ5ohMWl+U0QxG2jhWrlyqw5T0suhqef18q60bfq5x4VGv
jETL4zhIrDiPvJVpW8P4B5qixLkuxe9vd4t4ZscEr5FYqXW4D1wec1fh70AaJHQ1Jvbd0LCvxFrx
j2ySII2pov7X3giTkFEyjN6zlm1qOJ819bWGpoMRUSuJa0lFNG97yPhC3VTkAgy3gVAxzO1qvwTS
I0lvqc7X5h1F27p/eXALnzHfM5+MDqfEnv8fp+RlKFXeZ34tkMQowCYlV/1uiqk+/xPT3hPRtupM
+rhDBqzcpt1QIZGxe7XLG4cQcpcXzCj5WR47Zhk8NaQ2Bh8K4Lu/gAOMPo+A4e0o9SksDV13zkCA
m86UrU4JBZSB0UmWn0cvebu0uomyjSBC+JqwH1Nm5qhtt2DorQMrPJTZlZgy54NVjCiBq3PTOKUJ
UwjSykGG1LSHqLA7cWMUKBGQjGP8O3t8fByMOWI6JwO0lGADC09stqPndyON7blYgQKJ6PRSD688
b4e1r/dmCskpc63bE6EVEfnm0zVEEADQqVaztfyI5+hYnykedLWyMVNXiI9xFlslQI5fyx7WnAAo
yXJGkPYdKm8PVuqPTyDF1VaWR4RR0c3qgZw/GWdw9tr8J8Evm1psXB6OXVzaegrOsNuISDRrTvOU
0PHxvC6pvJO2Jn1G9fNNGveIurCRFkFJSwQPFnyZIIVloVLA/tf5U6PfRORqb2e8ZnKB0zZBJa43
ffIxE3qdKquDNF+bRDZBmoDy5zu5V8qiyyuGBhoI3iBcuoExmQ8wnW1A+Gdnr4FMdYWylvl+amyr
hnzUUw4CqX2JiSKjcvsZGlAnfDj2+XhIjTChZYyZe+HkQSJv7N4RmKBcEZhiAUFSEaH1L0Kxhf/2
pszcWL0pCFOkWSz6zzqqwjM69SS72rwNDfYf8oAVBv/vuJhUsktXq0o396zQps3Q++mT8jiSgvEQ
oM7gTzqj/6NPdpeNnwCld83by0so3of1WvwhV6vH+0a8bBu+41VfBz/qza9QFynOTu1U3BV054/2
vedRR1QdDLn4P1sZoYEVik85YoJz3SnxYEokrFdO1MU37LYOiLJ95ddxnZs51yRU0gv5arkqcs4r
hMy2z2ZcaBGIR8ab3cgsDmUHStTvInMbHsuaKauKOyTZl3mU9K5fAyieXaVeowvW1Q4eCSYZ/NEY
bycMs4i7rTNSo3YqW0AEVxalWQYEjyHF8KeCBc6f2ufYPFsM35y0xvnHMjhZWGI4tjibEF8yu3j0
aUlg/JKgGGwt8ofZxL1Fqv+JgyNSLqfcTs0V4XczDyKkBpImzIcX/gBOTWua6rd0DLMnFVk6u9Vs
mgyQPLLEUq/0G+3mgHs3meG47hL9OHS+eLE9dKjNuPFltDG7DL1d+wiFdiG5JY+PYu6Rpwrjt5Q2
xwnls5YV67ZMq/wBuOXgOsw/wjuafEzHwxCTMNWvi4s40IUz8/CMHfkt+aPq2FQ6cNcWZ1uZcqL8
/KpaNZhv996qiCkKEj7FUtuPTYN15fLKX8ocGpW3RZ4FhLXrPeRQ7n/f32aUFuH0TxkeRcAKXw/l
rBsae4b83El/mHbecOsz6fNfGAeDVMVUF3xbgYX1K5oglumxjycvRGZ4uK3b/YLXqN/ztAVdIKNG
Gy904luZbnaWCSLKvz6WtDmjR6+fd7ZKAGQp8DWMs+2DZG7hGPdCDAv+3qM1zAuLdr98okiRRmg9
YWsf0xo7SPvv3XYSBOzp4xu1rWLoFy6wu0IQfmKsArFCYzcX40vqaXNSF0ubd8MEA3GOpfWv8C1T
K0Gck/9gUKxVZvLztvH+3iDMbbAJ3N4JcWoHMYNQcZ+FkxoDV9n6K6ZMxPN1SxRhoJinM9wTK80F
temIwdh/zML8nE1Om3iD13QDwZl4syH/6gT6lqTBGreAeB8QVCq41F877z/pymqcBTgFG+2+mERT
B8w6Vr9qE3T3SUfRw7bkhqmogC3FabEguW+O3JUVU8QemG5ukzIo0YI6ZWO2Pu+YXxYQcScyYcs6
Ukat9GYBW+yljZtKK29GBGlgJmd8RvmJ6qsUh/wJ/j+RCL9lefblcKKUO84JjGS/ANrykyziuyHX
RY71nWpFjxI+bHRbZ0IVnK12PhQ6R5l03QgfnZrn1MM9XnJGG20cwbV3QBczK/pawi4LbGy31XX+
VXHuweFMdba8Wss39zk8qz9nU7Ze1iQjsPnwv0krXT0hxpUXrAP328PRKMMCBIHRsbA/uUoYS3sK
QBO/Z7zE/M8DcmWJiJSNPKviS+g1tXDeOEVexOCHsY0QHUGfopahW3FdZ1irD/ekTatMRvYcVir5
WStNw4QsSw8U+wll7Y281Uzamk9CzsMQyNAX8LvHTqpCqkLN4z0uNhDayONe1176N4a89Wtoh6s3
+yj7xKP3C7rF1rL54RCS/fyKOZQT8c9rXY31mltBF+ez/v3luhS7OcFrqVBxqT3GNwm+1wXJfhQY
6qebTU6aCsWYa1KCmuyjjFMTB7apY6bpr3RjKC0MWNkgyenpSLE86V/a9Fc+Od/mF+kvXbrEslRQ
msr54cOH9AIxbii/3XWTJncBfqeBKj4MonQIJq8OlgM3bKV0gzkmIablJ/fr/1kn5grwM9EtWHX/
7ZeFhzQmruBbwqhAaHXUomUvazZPI4nxIRrdCWvx7TLokQZS1k9B3sIYbWeK4VOux60uXQo9BkuB
JsB9PnUtswjRXRkD/ITqgEFJ6EF+21zofqLT4s0wQTPFtue92cLhCz7EWgvvxZdXEyYOaYrO0AvL
Ja33zXqrcBn/MCwzD9hOPA5TyOHqLCZEzp/FK7wr+lgGu7+cZDVdAIT0Bh8+su2Hdtel9rnfGcpc
+ZRNF1RpS9qJwPue/l6/YnaFjRBDiYxFBWRm+/Kf1SfhRu86C9bAi0An76iWuhs3xhuWY6zC++fy
glBgec5uUVjhql3Yf6FADYwSJhougTtMW6VPgVm2oDj0JkyqBwQZXvmi1bswn354zgAyxXTZumSw
mGiHa6yZ4KFLd67/Bz1eXT5bg9BzKjTNO3Q3LsU4SEneZnfrfiKp2GifqApk6P7YKH7Iaqo9hB/7
48ew/DXEPURKEvFmmIU68HZPthSuiaeQgX4pvVvCHKM+6ehq+QJOS2WSi+zyp3drJkUL2DHUIq2K
JnnUInHBIoxBYbE4GVDPoimVKzFL0lJu/B/RLDKGAKX0pPPCMpl9Thwd46Idavrh+cb7sZPpad4Z
pmKHX9Lr9vggEScrw7udnX8uftSc5ku0n6qhB9O6jpwPlTHTUy+BPWZvVG3HANW2/0KUwbouv0Rg
NO5LVDnVDvA7ZkC8UFxeibQ3j9ty8Ij1KaDr2neDukVexZZDnfk9KlyxOLviOrkB3Ht9fnZrsCsC
iNKOjHBpjM/6jfzDKuNEeToVZhzN6WZhh+vsKZepgMlkSmTAw3G/xsR2CepbM81CAVrWnO9bnZad
ZL0RTrx4lfiPgTzLezHvgmOPbcz37Khp3iJ1ka8bI9Cl3jFoGoPdArFHlbVc+uGy8zVut6Unu0qr
6iiRhPiw/psHZqmmuEs/gNHPJngucncn3Qo4wvci6r+MDG0IuzQTbNT+xadyP4l6lFMv1THsiROU
q9TK+b0I501f5RSNkDjGLzVYB9u3Cd4jzoYf0G0LY5dTiNbkKZlXXzqdkssgGxMBex4J0/NxTyWG
d3GZIcrJb4KIstk0uWAj6wxaaVKUcwmRTyT3+nDt4KzoX4JyZM6Zs2RWWWMILIU64SbgiY6VgW9R
79DM5k9rD/EU+qUTykO+N62OqvXPowQsfQuYbfOtsTvsdGwNz0DEYSoq8hhywIrsyaYUZSKgxYE1
BUYOggUbxhOhqmtKnTA9ZyndQaBYqa/5cZmFZMpb+x3KKvPptebVwRnXpJNO1rpJY+BfIQ91gadw
KY0UJDkuHxXdsQ8AguhX5By1RQcVWbE2U5g4S8mWZ3g9tUbgzyK7UMJNfxi1Lzx4LBe5yMamLSio
V0X4KGkIOqI2ezmigj8Y8FoH9e+S3VBxFyC4Y/zq/SqkD6vISpnfg2e/3TMAv3OQNGRTZhoQwV7a
5uDQ3drL7cA3LxG3qVziW+h+APxq/v1xToW7+W220hPrdYcAP/PO29+2eJtfPSkQwTYodO1ZZB01
V1MGezlDXVQl0SyVayIMY5mSzIpgTInVOOC9MDhtzQrtDGNoP3vKUtsefyfyMKz6+XwBYYjnlk30
jW6EnJ4yUUqvStkY+grJ9iHLQRKtYm2ntN/bPqb9a4d5Ln+sZIei9U6mrw7f8l3/QRvQ/a5XC5uv
+3q3ICxVad4VrTmwjMAxRHYg7NO3pp41AsXufTWx8+dagPmyBfgmyr2D8pNGHyOGFm9X0iLD9Dzy
O6PhoslVDzvyb7U69UMbHh1k+f0Q0L1TkI9FsTtM9s+hqg68NB4woFFRE7rcy/Q1P7MOzFPI9ppc
8Qw9BhrZwPzg+P0D82T5h+W854sOts20Y0dkT3CmDQTMstsuLjiXhYoiFHyCBDU/A5H9phfTEYuD
+dXyem/Kmq/U4j7SvmVx1K+ZbvvXMF4RUotmu/Gq8VUEbtaT4CtQcVUSVu9GQODFIVKL8WTiWJ+7
k7Gjory42MKK+LANCoHIQXyEXv3OObTtdLLOQZmcfsEDkX8iox+6TkbLdEoVCh3GSwqsRQSQekhW
J+5HYcLlNyRqbpHI4KuI8gpgiR5ISB+WgPPcJ6r+naCbHTdncKr80Q2qS11nnlCkd+AQ6/j0hZ+m
wSkB/TO7WzIhHWVt9boDAbZumglyGmvo1KCL1S4/OlpYe9fBEF0vvnN/6gShUO9mN5QEIrsp/eV3
AgtH34NBPo5q1QlvBzOG25lA1h7AeMQ/kcOtP971PKDreQohNeTD0NIe5RDPJ752HYoSlGuhoL1Y
v3Ot3xbAbgFCa1vQDIVinNyruwwhFqxc/nq2utcNV6CfBS4pm+v1Hyb8klJOTUqawaUR+QZk39SB
vDSM2CmOQq3nNsrWByuOk61oXkRp2DfkqfPHMQLZlSsd6Il8bYK/nUHE64EPySUBvqVMWGi17BEz
hxC+1H1eKd0vM9iL6fzKRgy8TCGGLhb30t0BKyQdgsIgo3PRFr8mP5+Rdcw5Dc+2z4LkDMK7vx8e
SGkfUFhPxfe//DrG7cbVr1wGHjha0JWlzy0W+w7IYXtnGGuV12Uk0IEKAjAzdga/KRzB0nIbyNFj
abSQjhAQ00Z74kdfsuf8x4l4um9oV4RYCnz/n+HZ6I7GUkJb4ZrrkdvVmQdCymX18wWYE6mrU5IM
WDFeIV4yJBAFKEAOtX/oTjG+/jdgonMimLraIXT3jEvvIgR8TBl1djEG0qEf/lwzX80dESfl658j
Dzq370NqHtljZLozL91Y6eiLJrr6JZBn84TCqP3FMb8A1c9Uv6wWrZV+ljkXzpRewxbo4WmEE0mT
KTDdk/ShJjtakCUjlNq/R/XXQ1OIJpmkDE/ArnPkyEk0zPweTQj75iB4r5XFn3SrjqAPpolRXavo
DRQqtZ3UQ/uEPBbK+u1dN4iziOkG5GZ79XtMQY2K8hU3K7bQ4xXH6DXiQARA30jgtNxR4pt7bZ+I
XOUcowxuT8QqtC06u1TmKrceVEi0dSvYpNCg0W69z0eNRgnV3/UAyC4vd4IxQ2QW4gTqgY4QEDCr
Mcd0jRIOgKcSZ0zx7Pnqjj3C2/MKPoZmeOx284tAPI75S4BNlcf9phEBr8EYS+AY4EvzaFqE4aIj
ygNOOCehM7dtT0I4XWVhOa6pM4eEzqvEkGAxUKo4/jtGQB6659dYBVXKkkGwAsqAcPp5iA4P3hGO
OPGBSQDK2Zwc/foUCS1+uUvI5mACvwdC823T0rGmDJj42DosshNPmEc+U55KHjBp0Z1aLtFEt7Lz
MCEdpIE5w5ptCiWRUvAi9KLDVswbNjIViKp5kxC85Jzwk4ByDq7pYnPFk2TtpVDzw7i2DExmwsem
TQRlup5vELo6w1N/VY4fAVliU1Ro5dl7dg638F/x8D7x3FTPxHH2aty66cBK0O6gh9+xCJCETg3+
jNJYyeve4Uhm8pDyBV7oPLMonySLDhgKQERKTRV1fLoa5pFzAc872MUEbXeBcTy3dGgG6UyleQcK
TwZGMcXmmmm9KG37cvRXQb5fcz6per4SjTgB5jGeaANzxsFwCjE3jDbxvTrDOsszYphk7hBihvaZ
V8qEl0dhi12cdoQJ/GmRbVKIFT2NhrMOlWYolFNiidzJHpjdagAmpJxxuKp9VR1xFvEzWjJ8rZtn
unCkOHvzFq9V2cPo5FEwbD1BPWyLJKgxiVNC8FA7nSlEU1jkz5eDjtEX8sQpHeyd4MnIAJDYKWyq
uka3r3mmIfQJ9737LouPIMTcvZoCSyYqPSi11WFdiEb33cjY6nUYnCr4ddPhXrRYNfIZD1stkJoe
w/P2LwIxkH40CCLc6ffyVJD8d/3eJ5HAkx5I7NeeZkFQyHKUh+VMumneVO6DBAsm4E1IUL3uq5T2
hegggIFRTXfqn/2JvGhT3Kv+XaDImiasP1Ab4J/HDvnB5uzYeukMFF+XEGBZUB6wqiYSlAsu07Ih
XuHP4iIO3jIdsGWAbM8LD3+L3MFl6Eb6KbypoQF+lEIDomXwNK2gGzEudiFYVZw5mKPGrTPDDBVh
byS40R6pKutGYGfnq+g2rI6uTQiTrRxCUEYEJRuQTqJ+oP7y3SvP84mCxS9Ox9AowMdhDtyXaOMm
94+xLGjI+5tVKxFYyv9S/yu6UQ/U0UB6bO5GpXaKwx2xYkynU+JyF3zfSXdlD5ONPIMlZzvYWdEC
cQTtqebSuzC7aWEzDWyrbX3B3bXvgdLizojJE5Fe81rFQ4jXfl5R6XuUBlZ9K6chVuBnOHKvJX4d
DEUZ4g+1ID+pZQRI/3vA+82FMvudzAJgj+90z8u8G+vRceAuIhBjxgfXg1KMobdq5zOEPzCEWYSb
twuL52ny5XKPjOLLZbvMOSMY6fpkQY5sKNR7FtR8HwDdT8OHyv2Huc/h3/CmLl8jPmFTaqnRXCTl
I2i7cgwUJ+Q6VFBPlmOyo3qS3SvmmMDWpCryf9pUYMW60gdq4m9RcxD/KEvgnFI5LO4i9VL2nHy8
+N8eU9vM2ka+oPlipBCS42MdDQGa1pi7zBajhOcOTKkGZ4dVBZGpqF702/hxhlrxsIhV5f5DJtbZ
PF8CkwRxiSBhhPKQ+KbZVQdmsMk44Lx5oXa18wLQJLKz979D7olJKfudKu3W67+mtRxu2DQI/Ohd
fyqk9V+651PZPS6CIOrD2oQ05+ufalcUEUR2DGvfp4UtO7vaGX4R6KD+eBtQCKQVoDcCeRnQ+W8n
hE2NsggDeSOB0qMShrrXAbGtuSmM85LsG5SeqioJDaDAqqBYzhnGIew9ZjiilYuG2nQYEiNgcp6y
Y0D2hUFUC199B0Kg9Z8hsecBSJng+AzJtV7WJ1AJ8TAVniRpr7XLp4YVLhp+BzoJ6pSRVywM8K3e
PGSZK8I/6S65lgAUbbCp8nrYy3Ko0hvVqKQOfjurHFaGl9cnYCNMSeS93wSF2ZGSCXLGE9FhBvPP
WQkZiwSCFSzIcBpdHhzLlWcelcRmjVsWWQBtzqdNVXIcGvw0oCfNm+O4SDkaSNfxssbBpCPHVYdZ
tVN7P7Knokzf6iayBreqIRWAgIfAIX1VxJbYL2vFz9hZ4esMWCYSAA0kKtNWpwfXerUXRhtvsdIW
6pKXcrexMHVZdwoE2grRegg/x96Yyg4REmvFvgEKB2lARryVqxVSf5FUAj1efqh+qUdO0khXgqaj
KMMrFPz/qbxEwFWq78u1pc1dCY8aANhPHnB3gYnMijsuYiIhxZBONjS3mA21tthN6d9Cnmuu6fqw
WtwVcJvIRBEfCRFFoK+4uuQJfhqunBYs7zrsYmdV82+fDc3HHNYzkZ2ZifacGCRDullCX4O++AK+
4HwHfrkRZOm9CrpRxTQkDr6joEZ68Wquq7D1e4BKOpzZSx3U2Q2av8yRNtfQnD4M09mBp2nLZmvi
hUEnV53LzYDUD6piyeIjODt2V76Kfxka7sHBTZGOVh+YfVb73St7Z0K7xMQOCVy+RD4CxqU0PmNI
AgcyKOWqeuA/ru95npmCEbjXunFg9hcs9cR+UMJE73y0h5O4pxoNigVFnjUSjT0x43mDT8B5xORr
rgr0P4j9u8FfF8/dU2ootzdgLqbyCsARodqhdxec98z+RGujnKUZH1kQrHDmt1PU7nwlnqx80tPw
ZSZhVzEEIKHxNiTKaK3Z2hYyK3AR0p2WpDO2uEJDRS/+DZk4usFiwlIaRrNY2Uqgnbvdv3ck0zAg
b2RDsXLrj+VsimCVLzOruqAH1SClI4CL7z559e2A2GjKH8I0GkpH4E/QR04xa7mMeK+QiKF6jFwb
/H6bVzCXoWDvB1SmMgdO8sW4egrU2oAvzMVzm6gyITKnhTfUuqWbpOOoLhJNuU/UNFoL+ZuUmXHi
ZHE2V3e3FIbf3VQiDD6TT8eh38H+snYdwK5Yd1dArraGig35v3r8yraW2k1rIpaYFDTBpPe7id03
/GB9BsTlwfNaPCSaw+lPvwXXu75oaoofx7N5A8Rq3Wu/d9hBV9AXGXQWSAOjIc9WD2//WaWsvcJD
GPmSeRKg74ABfPtfwMPcploKUqI/EjVgp6tasgdMJF+rKCBbzrOn9iYQcV9UDb2RDQdZW+DZrFzL
XJjcftLWssKAXAidGHQvSfeLXmIhiyjo8VF7vdOEe4ncXvahU8GHUvbLxJdulYvGlhpPsniCYwMR
Sr3N9shESQJFQatvwts456FLSEoqD1ttSSsl3bziqmjSqDIvtQBLXC42S+vLbdlDZtpMp2alhvsM
R+h8ozyxXWHnOkbmR8AjRd+4XnJRC7My6hahgGVkph3f76HW6yNQiDgX3S30y/SE9f04RA4mAW4a
9iVpKIDPaq1EG7vS8r5epYCx1UldvwT31BSysx7D7/yuKxvRWWYtqHsFeRDKA9k+bFKWGGTFgYiC
BnKLIOuGSQlbRWsPRsjOx1pmZ4i2YqJWOA7Y2Bd3gUQ24vbASTFfXeMqQqAx5KrvuWqLpkBdxJC3
4EvO71yHh2l4J5jBmWiPKzlEqQ1qmBkWoWEKRBwTPQTyR/qjDSEwG6zv/gad3nsFNjet0xZnMfSc
2gG5MUFFNULvHogdhopca4TUrG+yUS7ZsDjknCvYfjEqwMYiMT7FXfQmgIuVxxomxRUtQNpTr51n
xbjW7lyp+jpp3TQE5MjeKNeBlZE6ED3QkfFQ535/vDFVhmOaiiPwT1l6DKCKhmwDN6YN501xEiRt
qsxGsx4bbn1aGC0KxIFbCNVeMTczAPhXMlXQCSIrXdy2K2LqOVc7qyDD1g53DQPbCUH8jJPIBroR
oQ4FlS49A2NFq2flyqYDRf/dNvx+KFFwpnLKYZtmdEfA05FIjujuZ94bd2HeUyIz4wxt4nP2x/NR
D5X1/6e46YC/qAOk1F7wpAqNPdBh9o635jUCcKiCGMwjmG88gNGd9UWRFsKlV0nUjKTdka8zadA0
bS6YQRr6Z3xqb/zy7aR7robot0jsLkZzbm6wGqT9feXmNDiG6A/ZneZdF+851Z4xu2nCoUIs7HQE
frHpXr9PKAPyufWSssDn/GLKwX93DKXcCQXGrahaP4KrpMtnqYspAPi3t/7Qb8enaXBeK0h8qn/8
B4jPRiBKuYGGawWmOdPswEVQe5fkiODBGGpueD/LAvfDu+p47wec5wVzEW9NkwBqEJ6TFIS5qh9n
4npKNptNms726kRWXJMFjlO4O0tPju9YwhZePaxwApNGsgppmgdqFp1GKbd+SSwLm9CANcdoJlJ6
af5zQ6SiJohEynt/q7Fn2xI7oNwpHocHsS753pFaBJxeTUpTNwDMLxC90v1c1jHyRcoKNLyA5Hrk
tFrW0KBWHGUnukmLxWyFT9zvDIJSJDOzOjiHgxEARHgZGS5Bra2WPX9j94RJAFoMOb5IyEnmxW2+
RaihGFVn/MRa8BpZgZi/ofGS2pRQsOBue6ZjQRS0ECx4UYdqDpzV8Y6l1CLuYTEM7rRiB+UcsFqv
yW0DEZnEI0/BGLgkExZxg2XU3P4cdlrBJL3SUxJKHf2pWE0xzBuctRm045LX3QpNaZw6t09uEgIW
Tlj0aOWwIU/Ov3bsrzrB30l8MR03S9w40FzMiq55wPy+23rqvs+MM4mLky0jiUeVU3+ypv0TFuo1
OGM7afw/MOwcTdXbcKjixEKTnJEzCSp7/7WsGXF/n9vAiS76+HsUEaOWK8N6LZATGilO1Nh2X8WG
iRipsM4fjTr/r3zEVpp8CqqjBd0Cei5S9GTue+19q1PsMrWlTmBLpc6xXFpqF2fCrJHjVNBcezCu
+s6p56pe7FnlpGXFGGtJJOmQ9NMSuSITbGerWDUnbvsquNYNskBDEoiau7rP4Z22tpapy8IWG/v/
z9sRViK7diE7wsI1JwLcrxbUk1ImASkj9VSj1ynIHmPkWDiNt1VPnDe7DoCDeuVywHki0tJR+T//
nSVID/xFEl4/xMQCagsF5rvScV/K1olkdKoFsK0It/CV1KDEQunF7mYwWsAnuP39C+cp2WyChLHt
TarIsRBtvHaad5I+9qRkBqNsSQWwF2b8Uz1iPflTxMYNciaa0l1+PHyMPsEfDhtcWfb0Q4QO4KPj
XsBTRXFzvqOiEg9sUCBvbTzxNfMQAqcWBsuyg1J8TTpG+4/UTMAWfvY8iiJU8mwk4ReLfKP+CY9u
vZndwwODzhKiNFPtkWJ7yImKJ30MdwZof4hUE+st1qE85Jxn6ae+/AsvW3ZcK3co2dEvJgejT+Ud
nrBP6xAlyUCKWNtGG4Allm4yvT20QpVE/nzdO5VUOpVFwYg61Z3WLQJDfymY/C5IvuRk6sD6n+KQ
RQYCAOa7lwjxaixoNuO8O2SFsOz+5xjBeNYDqlVVePw6I1Hq66sHDqE0Q3b0AHTom9SgncmtIpis
fWwx6KQUTdi5Y+a8Yl0H7Ypuwts4Pc1QoJSIcnMQBq7L2n6UxpXuLl0DQhcXrEuU/CO9mgrnVzP1
l2dFeEuqi9W2YvFJbq5GOAJ/OZhPVyPe7E/L04kTnflgyH6yqWWsAW7f7ol/s0Uo8JsyRcOq+Pke
Hi8m3dEySZis2W6gGEqqTzF4rbVB20Rb2YdHgxXJifXKeP+6xvUH/+vTjGo6Uu1WhBIEPqUzF/Ux
Xz4HDmezrQixNT5O7rLVQ3uHLP2TEBxJP6TEHc7Xdm1He6sYj4JZ0LAj+SyO9/nvLUhick6MPiAW
FbTW/IUBZItmU+H1spcW7oHhDmiWbj7cNB6jCnxQj/rQzxiX9WDdgwvW88IWaQi4+tVHB2fnfk3N
xU1vnZeASmBVzHnU6MVTMqAy4sg06SpyjDLotLxq/Igkm2IM1Dw2+EvLnsBwtg4uoOsZJtaryCpk
Pvu0xJe0YAOxzupYcRAQM+hUXmJqnhwwKcE5WnnDmP9L61pE0z5f7frBaM5oMbMHH+p/oXcu/uN4
kq3gGxRw4ITmKWyzwWdpecZg87e3hJxSC0XTO3++kC26AYfhQg9XTjhD69a5wF/9ZEAy4yYb7m+E
AhAYV3r9vezI3Squ/7ob9zgqXf4HFyYcUCMwnYEzIsyzDpHZCrUvF4CecDWcv5KJCCoPzXYh1Gta
6HoEEnKoOj1OzTW1v6L4XpYaYuv30QFC0Kvedawc6Qa8mD0gQsODNZtriq7s7n83u4qWJFEatFxj
OZ/zmmE8CXmbSOPNgSEEX4G6YCKKLgWY0lVuQACWN8fyPJpk4547wAxAC43xyCS4nR1z3u46fA/j
QE2Fv+yKKoK5/0JkRos6guTSM4X7O+ISsyKaBjDxGaYM9kvyRegPr1IJqlqTpi97tC4ywTFC5xha
96PLB2TtfXC5YEJt+HVA4F3FLD3Y9fcNiTx7EZ9wwbeckXn8fr/jqJOkyZW/wu6WQNYVWxUTqBIo
mt/vMKdL7LRSDDN2U+8XclkLY1OZeYhksih9sYE24m6R73bI8dtP61knCHw3de1mx87RQUSj8pDi
ap7tnrL6sA/HZh5kkAm7ZwgVDci+utlJ4KFUohWuIDzTZN3oWIvvwJF0TTtSO7elLQnwGWlEvR7t
1Uai34+0XE7uXJRXgtoNiclfAx4VOVjj5AoY1GPztn8JxytxQ3tceZwRwAwoQ5YU42cbJoUOTxHW
XCej0RDtG6GxqODhWWIQFvGcTnYvlGDYbOxVp2R39/i98ONg25nLCR2qv1m4/BKeI3C7YVzCPXbS
1uO5KP67015JWucNxhCmMOrXGCjRfmyBTpOc4Uvjpx6/oFfjbbIHhZfNzLJuywfIGWwDjyXNYwTy
32JfZDNjPGY4lF3itHtT5t9zAjRyvb2riP04FAPRv4SmodibUP4tauup4K5EPjyaI6dVSpRWT0LK
G3TJJhqOe8c4eexglRR1UcoAg/Nm/oy/02PQJPO4xCZFVCVK/QnBO5hX/llXosKFoy1ZhJHmA3Vx
r6q9Pb2kF/vGU8jXANCIoA4aysDRGlj0W9Vc3zZBZVdsKrrDPHa28epPxyNHmpAUbS6k0eqmlvtA
qmfoopjulRz8dHbasmF+2jwIkAdaex3eTwT4IcVzd4SrO1pt88ik9XzV7UWaA1iAk+PVzQRJmwOU
exWeKTYuRVJR+VBeqzYftMGiqL3HotATEtw8tk+ZipH11KZFHNwSNUfbKdJ28ag5bVmOdVh2mdAB
z7B94nXDJCdpbBP8t4T64Gz689vQmtUcdBqB4V4yfLkcYR+4FpiXxWmDBNRGTd9Tb9WRivJc6tpP
+4RKElMLkB+Uv9ML9YbTavaBESC1XBCi3QK79lsEBI4vGRe9rD+5f4HFEcfLeapWhO4XPi/RvbZ0
NKNwfXadj0+HeEsu9JmKFe9TbhNkQJq40LNQ42dkBwYUdYB+1e+RwtjS/JigwMm6xNuQ4zX9uZV2
XFb3hxmllsaMCFR4ZgXbpa+UnTIFQafv6atVlu5GeiKB/N3n8a7Pg/Mj/d6Tn/1IdmesaX71sVpG
0AwO9zv2c9bpJBrnDPzq3+BUZeIhsUM5s6Qw0WTFPZMxPGrb+v0S8kgoHkYbryxYhtE6xJzeQQ+2
rwnwtyRL8MDM0RT/7mm6HlCn2B405hA0RdmYe59b4lc96ffEO6C6iCPfMmWyfgpGU8bGNDjxA3b8
rVrQSG61UwfdHERSAeYllxXap9of5k0KP8QmkAxjnmL6USJkrUnb1Oa5JQYLPwfyikMBTlIcz49k
sDAhK5GGuYGfkR4Jacb0aLA26iEbA9pxIgS6y5iExpGbbsXSF9w8z0qETvf1yd4jMvdcAD4iP1hJ
tD2Fuq7xYbqGK7vuq6nLS26LUFM/vh2imS+HgqAQG74PXE+56SuIRfLZB2wQ/h/WEO1n9FVtFKYR
F1O81sR4kuYmqqGMv0RVu3ya1Hktgr+Fic1ToZdFeR9bqGH27qBGe0QizLlLTjyVWkhDw7FWTQH+
3lCHRmlcORVSuBCazLfH48JMCxOGrkLI5gsdIaRuouWA+Q3wmVzcPPS0W1hIetbNjBzFZT7QBj8N
wQJboNDYOpda61uqlSeJ7Xd5kCLUBOT8P47+WQFQuNZsNVMCSESD0qN4NrqC0E4qThKKereGWHoY
xdHwMecW0Fps/QEAqKzaYH6EAURi1LF7rNBxT1Ebhp6GPa4v83/F2w8hu3BLreL745r++hIkR934
nW1hJTnlcGARJx+CgeztQrc7q2cQkVZ2y4VS1duvGIyUaY0RFJtlau256XSvDQBLFbX1ul9EZS+A
7cF7RKJrv+aiYLOXvzmJZ16CgUEQfAwZ6r4q6VVZktKNNy6ESc2lh52IX7L7QFSMQeWUCqyp5861
N8f0J3voDZxwj38WHhgirT34yC0FqfRt2/fLr3+QCRxADG/glJyWmPTeL0e4rCfFvc7ooBHTU/HX
rtS7sKLFzZQRSWNmzfc1HzMz3wPnoOgD6Roc5k1soCswCo2T+NVEtEYo2L14C4nZhJRIGnK+9ZLO
jUu5qfZWaKYNA+rOIVR2QgFrKlLWXuiftZF1sWv4U6ENIHmvFZiCdslfxgnjMQyNY8rzg9YlWvek
lBamNN4FSVb8yoaG36Lwusv4/hr3NNIbgtfgATS74DuxqFKoupS1VHPk23ZvDNS9B8qdWtU4JqdX
D0atxSBQCOmEjTGTVcEnnJCc/LSVsdIr8RFb9/7UUoHD9f8mkcxNVFyfwvot/ffek/G0A/HfSn1Q
2brdFqOuvNq4e85nuAh4DpnDRuhl6WYDfaPN3ebimquliNAFnRBGymKeglteMCNhXFPkvx/LsAhE
g8NCdhHf0orjK4mLuNe5C8y4Russle2H0qWfE4GYg1APqhH9Bfw4a5v+xysU6zLz1DO2u73dz9ij
psvYwDpjKxtvpHqgBApY/6yLA7yn75Z2zRNMBS8ccW1j3yYAKqb2Y6T5ke2CE59jFDL8Kig0Zbgw
+9zZiwjaH9nwCFuxiPH5jQu35aW6GXS+F/y5ICvnZ+gpHzdUdKs6bCxJtZiIcXSbo+4fKzuyusgQ
rmDdsCv38+/Feab0dwhrCzeKYXzfOrm8FUPLLwBQSQ767frPTmPuTqH2AIdtmYdwihvA2i3Fg3gy
CIT2aBLicCwfG+qm+HMG/p9Oy0nEOy3RbBhUef/gmLWgLD4FxVocyuEAA7dXhmc+AbUJ23JvxUYO
QYgfIrZAoGw5XaayRXGs9Np5s6PygPgvgTMWTR9OjO/zbk6/Fd0N692EklpCNNMHems5RQV2hb6k
Q0P8SFL70MyeD1eT/6EWvkPhk+6e2oIc2jrmG5rmZJvhG1jDj5W4No2x9cExyBehlVQ8ZazcnIWd
MPFG74M6dZuyL0AX1pzcEAaAipeZPUVXbPI3D+wTnODiiyUyv8ZioweMaViuZB673jZGLjfrGpHi
iHKRcqbD9xy0MrHtHTWkp06Nf/Enq1zrK7hJSFpzPiXVZ617X8wm5Q5lzNoWk0Bbpvi4brPGqA+g
Vw7Ru7kkkml32LBWUoVv2ol7O2tky+0F3FM211Ol/hBceTdHqJlFi38Pssebnr5z7EgkXPgq45be
0ZCGbReBuWKWLEaST7f9Pfldq0Cm5y/UnuKujoLbr/gVwuG7K5ttAKD8N0m1dvfNosBiYPH6MPpO
M2s0A6M7gy9kjajJe3JfiRes+c6ToaR7B9ehDOEbwMkyOIhG2Qm3//t56CgLaIev2FGYfyE7LRW3
qQwQsivltujZNCknqS78Zi5s2WUapcXAD80u2zVKeAhHsGguZ+yv8WTFDDWHAhYQ66d6X8JDM7HF
Lt+159N0nFKgfxA26DjLw6hEIBIfZbM0jXzuXCYF7+XkJnmrgRd8m2yaG3PESkAEExEyPmIZN/ZQ
0qtgYE/Qk8IMWZMDqqSiMI2EVsNRQGA8+UufMyNKWM0uCN6PDFNoCWrlzbkhmiUyAIfnlcrG3Y+b
I+RiMq6cxKeoBMJMk0ESctQEEx4YM+CLBYo2+Y9VvwW4rFNUNJxKBjRdMFz3HLpDnCq+nhHhN5TI
hCIPM1wumKqSu9EGCNCiKHH3XUHnzaHxatmjWtsT6d0CwRrPCaS+X14D5xEq1D8h6aYV3vkBkG1B
qN5KZ0CREMYiHPfjD+QdQP8B5XLFAOzWKp/WL7XALUojE3HQeDU9rWItFsPR1CGZgXWGCHlt4MG2
aAYIq9w1QUBAFvjQlBk6GeyCrahwzbDZVb3mR2a3j8qtJpY5zh+R22G/8AtgWTq21A6aNT4t9xbv
WUaZyEJzL7w83ma/DEQnl/NOY4YjmMi3hbg1FJ+BOTJytbBA9wQdQvGh/d9/UPiix4RUk5esOW7K
uq/6mZqr+HyTd8UeOVzXb42XuHE3LabYWn1x9lSsDwG3iH0tIvAJAEbSC0CnwKl4Zrv97J1b20l9
IKWFCKDc1No4tFCsBAfhf0kD5obfzhL7Iu0W2nmjNkZokshjL5D0xX1yW4TzVF84Disi2l3Yhs3o
0z8RPmsmgv/wgdSoJGoKnni754FJnA21WKqlyFOdQEz91Yc1+d/SqduDhydHZPDNnDsD1TFJ9ovr
UITEgUzdlO8LkLbMsIL/o70MU9Y2ca0MwZWJC8Fpi+4q8Rw++VIljTcbXbynjfdFLDOgXye/Md8R
3PxDpojigIxGHK7mg7kRjme5PLRHMAO5VW6S8NNrlEgHhVGZte65LIkWkmg6Gia0XLkXZHdQi/g6
qimAZVlnZ4ToviQwdMF0CHq312Dlsc1aq824XngymvLqablFa0Uy+8u75KVnFsq8YTL8gS+rqRc/
10gfYam+VhBOM+Xy7WCH20G90KfqPVF1iCrKGVSkcZl/eCl7KmeNUrkVgVABo2LzK2dminUNstCM
+cK918i1KhII3xgOJmmCqX0DSzniQVVD/f9s6ms2kerBhtfArl2da41Nyg71pMJPpVcP8jxdAesv
e/IZcpswYYOKlSRfj/RFX05PoxNJ1YQOkK8d+B6DMrIjMFX2H4GPY18Z/tqFbb1eZ9QXd+6frSJQ
BzAUqR4FjUlyIEkUWZtBNwjx432sqT9EkDN8WuliyHj2FSQ5hX+cXCzNa2Xs4n66UkpOHtoLv/z6
BVxltKQopeGFtRboIdU7o3V3LNFlJMWDJ0riSFQhASt4Ximsb3u0ZyeOVKHpCjEBdwDoFzSO+yKv
Xuj+kbz0ZlIHy1MhJWs9V7qy3SEXn3oEfh9ND6JJEbn4mIwsahulUZUeAKQ/LxrUlTJU5LPjNoxl
i37uQ2mC6zOO1UCWtTVYq6Fqjot7jz/umbmh3/DM397+fGFYKN3jaP4UDgUFhfxmRGMEuo427JVf
yItdaU/1s5DnZPiY/MuJErdIWWMd6iKptonpn/Wh2zh2lpMqMNYnpIOjjqv/w/4hhjzbUjtc0rMb
tqHTJ98wKvt9HhoPb5NR7dI0YTspS0tiBDQ5Ce1+8cd/wM65T6emQ7hgRtTTaoVnsMeaIJnwj4hD
KDzJRskwA1FlwAd+Qoqn644kXw+7UgqW03AdNXFnpsGzqZ9zw3J2hrq19EYnlJhjKiurA4de+FDg
Fpc1WtcUDWsT36RZgLzCB/r0kJERbJcbY0NYrNawxxn494SO8DyKjZF5sAAmpkLCQaq9BACuFRGk
f7+gLmK4KWNwXCYnjnDM/tCTKzNMrrKyxG+2eJL6pBLZEKKtB1SkKJQaEB7pUUQSPbP7xyiiNgwf
h+1ln/SDS+5z8RQ0+hQ1dW3g9xKM+hpcYc/i3BQjTJOBi7kCAcXjoDvY5icGEW7JDFYHW2TV5LJH
DH5MS711ofE8DZu7Gl6i6hEwV2AR0POiM2NqJVAqDDCg2AvPDWyvyN3EKMs0wxZMCMAPU/A22scb
qK9jmy29z2S9dw69RVoOHLJAHz0ePvfXY8rDfxVUamOfvTtWvH4cwQsnACjcDF7ZCE19oYV/LtIN
fmbO/jOPwk9K3ejanUqbAOKa6UxJD23tkJ2E2iIxhhvSXR4qzIrbNlPv9RQPZ96nPJPoPKV4SrnV
2+HMunRM+R1w5+6OjYa5uhaoD10EfGT2oOfj0ieg67vprLrbUiAWTxTnF4tZ31RolMpkEqQKDSI5
iptHHYipa0x/G0oaKn7RBO771WmvrtIs8JiVo1EsuxV8VLraQookSDTNsmfK6dQ+j7oZUj9eFnP/
FRfbDvmZ6s1C2lNBYr96Tvsr6KhZ2p2GpgC2e3rSE+6egEwYYYpVlaB3f2FC3k+UBi561lq+ve/e
wv6RxSlApAB7MQVTUhLKvbwNwqPjNOfz4hUty93hjT3TsAkHQUT+Rtnkm/yPkY42WdRfJZMI7qlF
1ch0h/GEucfG1cbQ86EugOO/CqSYh9duDGfDu4UKwGdtelcUZa0la3hgLJ13J2PsQT8YCLNix5sh
G0XuTI84eAownji297OFg3bQV4NqSadaSGQnRfP2uFjz6rcIg75WcCMdIIxQYSFeMTz2CmXWkS8B
bi3fsjc0dL8U8OycXgqoGlcOanfR5Bx1W+mTBN1iw762fTgC++uChjTdQXAWOdHYbqSRFMFSf6HR
zP29cj85SjNX/WfCu0E+AUyKXNieZNlz/cNdW8u/s2LITrJnc1nTBCPsczFb/SV8Da/y92xJ2kfw
SGBKjGQfqtT4QYCRFixAZii9vu0TydWZUGIvtrOwKIFlfV0GR08+CN/z/iEDn6gQKMkM7yfwDrqR
ieMrBr8DvaIMSabjsn5R2sLuovrA6RZoXjj+zg+LWbExRyiUnWLYNa1G3cvofLT+J09EMjVmzLDs
QLt+OLndW7/4Zgwpnqx/4X2wNCeZU5MGwgtrzH0sAvTqmEd1lFlWo07ljLijkV9NQ4t2Z8Hky0Xt
XeUqmQSkw1uc7jOm0WUc+wB13x3WC3wl0nK5liCD11mJgmYkKWSEqtwor214565Fx02qjuLtBv11
2Q/s+R3x43BjGcmCO6gPjgCYhz0kibbUcR1dInWA4w+ILWtXavzXa+kArKc+D/NQsot1FcdRIoJq
iSfitYOIvIj9e1VZ/cWxCU5pzMKPJdU7wfDMrYdzDz02dAuP1j2v2lFQdp9F4URKnznKyTwtUs+6
CzqGZySPl1lCMjGjp4aOZD600tyrS9wYNv+hSI5bSL+vEQKpeU315iTYADkUZbt8wMGsMHin9jQ+
p6spL+m5/aN6BrvUXoFcVd0HCI2k3dZb4yi/LkKCxGcy9k8/p4Q+h61yx7/5PtaHd2+NDJ1km0WZ
7kLTh75XIMadhREuwvixnpmofkiSj8j0zFVWin5/WtCQ/NT15VTnXg27vRfXqOb6FQeIaEm2RpKK
NpweYVS8O7SE+ERWTQfTly74yAYNAOpMg7XX5S0kgs+R+YKW77019JvasNIJiHSW0lxAHZ2x0kJr
plYBVHq2dMJMPK5s9soInzKjj9iTk+gQt73mDxIix4nxIJqGhTIh5qhWToDnMQ8hOoYUAxz7pZLH
6LmqRu3EadgTgqR7+Xw/0tkGTVd/1Upi8Vd951UJKVJVP4IxK68Oube0i2xfUhif1tQ6uXs98gTE
g8cm8WKrAB7fY+VxszSxqSSamcnK7XF/oBdZ0XId+N1V1kvJxu4vEo62aiMB0ASrFh14RML5wyth
0Xw4Nvs5YDaGtDvgO24JikDIZvPnePQ4EftA3YvTNOWHRqIsbfN3CR6ew5sqNETEp3gySl3ZwA0o
N5PiZcaEWWunoYx+OkNaZ+udcHYtbUyP3VLGi2rT8GhD+UwNTqncFS9/vt2N4d1khZJ19SYGqh7L
nzRQgpVS2K9U7vprgvHEUAgbSVMKsLmMG6TuqTZS0rmO3HGY/rPmgscUXfidfTH55YQORc6gUEm+
Ne5gMQNKxYG+hEMVUVlcHw0QfyRK1JW7VS/fQ8Uqc6MhwID8tEl1ccN2MM2Eppv9KEicC1u76kEY
cHPCjPyFmI0q8vdsFpC8Cd0Jylq6Yu8U7y/GLDrBz6KSKAtZa/NQQjIhpAC+jutRMwFq9OB9yDQl
1dqsqUKkuO+SiJZpUwM8pxW5bwUBpv9d/XtFL+EejLopx+tqkihcVEiHgPcuZxxOU6ebCAdI2FgO
afovDc4ddpOk4AWgq+YAG9lKTBCzM1GgOti9rdRbxWNLHDtngdTq59sC5bryGMmYzwjFQ99Vjs0T
qMLeDGwymi2Fo4BDS6HdGlJo+SrTMTJAgGM96QS38bMUiy+rgP/bwLzEQj95Jl9UhSRfUOViRSVK
8cZLO22s8eAX9xC1iyRQHyaddK0tW2uRiNagPh/iUzmyzUVcI/JXfgm+WU6yTOUkGJCU0WKblfNp
lQ9wAFlueyNY8wN2HYtObb9EjweBuGJqjNIl8TN1TG8+TCLxiJhqnnIpkYSbBpyRrb2WUeqz6kf/
LfQ8d8Zd2yBdBBLkKkGHA+jtSKP96ue0oF1gemEScj0Bbm5NHAN2VfDWoISveY4VkuhNIggi/HR8
V5Nh8QsT+cZvy7IqjceSW7ou7WnNb8Q9vNdaZRqwuPtssX6Miz3507uLKHNkHjxVCKXozGrPtBEe
mx8RnymjHTNtDY4wyfpLyoK8VgwacqTyDWNlc4qfKmnUTz6QZkJlybC8xY8ozPNB7B+SB5cOQKsA
oyNaHgFE1Ab+2m+AGta5KPsA7rqlHry5dQjyC1WkBHoqbgiGwCwkQmXJk4ehkXj1OYFPjz6HjscI
J0nonUZaEkGBHa/mfESULkPSpM+CoQ2mZmWM0d+eV/sGasOiKWBUVj8YxcR4pgsE1sixB89++Rt2
LtfJlpDMRUigvUKBOqrdAHdxjUc0a/jYo/g+05lo/qLkDmUkTM+VNCGpXJ9+VSy2RzFVanPGLvTB
v/GqFsRvjzDdWc+EO0v9uKv8gLP4M6fVgSZAnBqMy7V0etfzVMET2b2J6emjyoLZp4q9pvwtbXtY
fli2jZ4IYEc2+E92SDdeR4oU+CWHiyDbHPgeKqYK+15NwvPwJfkP9I0BJmEUWh4B9umyk5qwqK9D
GxdF0Z5HYR/1LH+DAFFhAzxIk3kRJw/z6rnLq5F/w2IySvkLa0n/BuwM7KQoNWiChF1Q8Q8s6+/7
l2AFk+RPbW+OKoy/IlQfKPPRjjdxYpfOj1DLj6H+zm7nXrKY7/8b0O9XVNArnGtiPymHlDpzeafS
E5GlZkCm2hncxUkAojgo910fQrbyIYVQEMHpT/T9/UITSS2200PBKQgGNs70k2+/SeTbvQWjS62y
kl2i33tYxUkCIASNdbxGbBtfAwJ20iN8z9YMvCuoC/iPQm3fDEo1xh0fHBnCMSNI01o8WptyIEVE
UBD6PBiBO1YhxUjHP/lc/nT4snYMYdihDv6QH8Xo/VBFtQ39pKpCnPF1VZdXSBnMn/XYKqeaU+9G
OqYjSTCf5zvcR44Y//JwzsbzZWALy93rju7GqpQ71Tx5nPLjMlvyuQ8yBlJA+9kL5ksuoLgc3S5l
hlfv/Yix4PG8oFaAfdekyDGmuMblubi4cJ4tDwRYRv6+FcaO+rblmqpMYR6mFgByrztznPo+JtMN
+HO39WPc61+6A1cWPMe6sl8YDfceWu2vjmTVPFW/kgzssbOP7/YFXEvDqs2twJi4uwcOn9lPUFaG
DG2KjgssG8dCI1nyiZboG7ck0miou5t++/1DNHR7YstTcjtHMWLceEgLHqB5AnJVHno/rkh9iOGw
WEqhKFDFQWmwjzJyrUr3TlEJRn8LtWXjEDqG5ZiotEFLqTcKC/XJL6KJz4ooLdZckGSoi999NJ0p
GtsQa81dY4T/CaMPC2NEXfVoYPfEuQCD+ALhCZB7Qr/Et3axvS11Gw3LDU3ANaiu98AzJv9ZPdHe
IDKlFrzbDuEVV8RBdy9gesghBPUOvP9/U0t4WuHHTra5kzMKYkFM6UGmoOmUqtzUH9v+xk3Uygo7
TZdCt24OqIlUPmrhsKg+9mldarCY6LV4sqGxd07fXELDxTlA4xucLFiPvGnpH0A5ZCHFy8+aBdNj
qG8sYSWLYPx8j0Lz1G/vkaYRBuTkTWaHa8yuqMhhU17znYnRFhpvEY8oxJuaNLDXx4bdpmICOgLp
jA8XpXQA4b4x2ABzr2e45U91WiiYPcbA/L4F8vATvjG4cYQsn85j0/KLJOqaEnwjpXzKbFt5gxJr
hOC87C4DxS+nIer6uxboz57mr0XYL1Gw3+x3xfJU8jQVvNezZ0g8aPg127l7Z4dNINJ79fZzfpQy
yLgfCH2lBrMWPXsQcTQLayWZfBKeSFQ88ZUpAAI40G87SgsI6qwyNEBCbWoqNFTs5PNdn/0umNt4
yexvyX+TV6jK/4kiloT95V9VQTCfQLUmCyGGktAIXGN7sL4ZZoIRXI5L/05PkKfr10A5CTfy4D9s
pGxPOIYVhE62e/2USXlNQORArAl2kWRGc5I26RfuxVMvSf8e4HIUbVKawDL9D56EPmhVjMl+nUTy
tfgzOtADRxj9BCMbK0nc2UaAmtBdxen1JzaM2RJYMRwqnsAI5a4vJWDQRgu9wJQg0zMlRbnOzjjM
yFqweVG1SMiSHPV6L8hVgf0647ojbBcZ7RjqJ+kosmXFAK0JWEAAkUN6LdDDckzrorFH2kCSDNWM
vzKuYuXZ6Fv7RBo8zuWT5OznUXsSQFnZZl1fd9edszt6yKAZK0BL52BcmOBfBewLSeoC5uyVTI/J
whihvZbJEvXqUpk87CqbGokkDqNQmtazhVmtmM/UhDYz/UX0fE/uzng5O7KvdWYvG+8vxtbj/SXq
+RcVVe90Jj5/ibAJepSEsEfq83CFy+TjI07fPhPqTDhY/UrTVlT4IOO1qEBFAwiqWAwJ+FYb/l3+
ro6NU5b9YgyCl657zl/kBlJYupQsLExjo/PomQN2pjW6fZKv69vTfAsX/barhcZ8MjkQIXciv+Dl
e0Fvp2zj0Y1eSP87cM+Vw9zAVThqb9f7/hKNGf7F1aM9zNodeVSrabt3KUeIuXBqDAi4KZI+vok8
UcnY7yrOqILMXfZiedfR2j5XqBMpwa5pLxNhgNj3j0IfBCkrM1PyWcZ8Dq0fYvEX/K0bbeYHmr3B
RHZ6W6C+fE9sIFxLMT133P8yT4XVS5vL1+Iv6fZbG0CfTQAq4gWtpQ8rse+qkh8Ngj+IrAhBsuUu
XMDrPt9eDCyYWKB8b0A4ORvON3i8POPc2zYCfNa4D/VYlr/r+QQse+cGLSJ+1TvqNgZuOeuj9VvZ
N3G9QQjxxaAODe4CqYAT+GneFAY2398ba91RUkua/G1vQbaD9yJbh1oW7tmLsk2+yajnZETyrqGb
Hj4tQjRuimDk0ZPW8jsjl+hvISnKPcqBSBe1UdsOcw6gTYmoZnp81+kk7J4vYCoYPlyzrb3JMV2k
LRbDbuO0vZeMWfc06ClbcD49cRZelrAvjhiQxAI3zoiT4PkBxMRUJ6jkgPn63oIhJtuLRAAaUDep
nNtNMq+H3M6pVP5s7D05k+a15lZNd6J1/UIH1Dnb0b9CVCuMWAbw5DlPMBlBsa4BRGuVQgzxkN65
OO7vw4C+8qyZOrtHqsuzc7Y9ex2nWmbuyoj/R1bhquVd1e9fMgpmXzB9fVDpb2wPD1OhRU62wusU
BswoNocd1i5340J3+IgC0U+MveKSVvizI7gOVk16cIxDHfayvAyt7T0ZCQqsQezA1CKyTsr81lLd
l2xekfrF+thboljiWY1WnqndRimGi14szEIGUXiHOBmUHZGgS2DkoxuJw9J3t6R/OjE3BZnmhWVJ
jehqpxBk+qHHiVnybUwhlXD542Fu+ew0oe1Tvc4T4LfbIAZPOonlvOCdzDzz6QSys60WK3+sZ7Hq
SRiJTn91ZUjTosapav2LCldCHGKr2SPlsn0HYkJkri8ilYAVxhOImdKZP+gxyKvazDGZQGYNotx+
ZamXq6WNAY6+jRrwvU40S6XcvjyHHTpDLHUDnwHKhyC0/xQUAAZYH0Lx9U4jMGmFpXbYfyKN+8ug
8iEnuW3XDoyFbtHQXqtoPPDb72Vz1JoysRsTqPgwYAV5uCg86aR4US7Xo28MfTmxVtJfpo2PsOrk
4UiWNLUPt7x8/tZws4KmJx4bF1+NghVSplHl1jWlve9VXW+hRiRV+i9T2ptLLSMdit+1dzPZlMhk
SbFt4WBCLTAt3Vg+qmF/2PAosxlWHRrIEmzvP8BKJCRqfq7Cr/TuRyvQfrD+eSYi8tJcTuPhvnpT
X0TooJ9OZvnS4oC1taM5A5ORT9fB26Rv/n6QHGLR9lmlu4ZNooq2WaT6zn6W/Qf0QsAZrVOE/Wnf
Qj6NLnYbZ7+DoK0OetOKrEbCYNSMAdE9ksgDXd+uuZSZr0I3surLvWbWzyn6M/j+1snG1HotN7cl
KY7dkkpm4FWy8ZUAAebktosMpzOAECR3INALFRpwPKascAr/MHZfAmCS2m6VWt/tSMPC0juvZjyR
vFf6CvkAawwzHXVsd2KZHIa/Rj9dK8WhYTAIHcfkS+ut60eSth1Br3yqqcYiMuRyT10YIt2SLOC3
/JoO1+4QdT/k1zant3SPlHjMUWRecFHdLURK8wCwTtNaT5b53Z4KtrY2SJFv/7/1yW5Eu5EaP6dY
pwHO2ESNH0SWa3Ziic6904JdmL8YThxW6lP2AQ/aoYO1zB46+u8FtoNKzWr4/7SxFon8DOpkTlSc
CUOiG8FSACxgwnEx1MqlRlMzRHN6kSEGatAiyGJj/PNehPxOVlB0bYZi7+SDXtnTytP6aMK32Xty
Czi5rhsQnHZLFTif1QEoz8q+k+/eEl1rcMoDKGfNgteD+Eu8gqw83E/z0JbfeO7ZqwpxGVnMncHK
wlxGedWAHJ9X7gLzFEkjTebo/Q23FEqjy/ccET2kSDaGC8ZxLK99cH4WADisF0kHkcWYJCJDF+wV
2oqWQwgzvWFIx0hT808Xi1mKIF9CzAE1JMA51tP2vs+Pn074oBuqGNmJL2mgJT9Nd3wQWgaA0a60
md7E2VZWidX2p+pDWgg2n3YUnpeFx1zGhLyaEpujbYiu8CpEBI/2YJcltqqalBnT7i0Fv1X4P7E3
NUe9NXObbN1AW2l4WlTWXQ9zw8ZMAVC7LmZZp9O8Fwp0oa18oCrbcAufO1kdPCaJ42REoZQRQjoe
/4Ex91ZWtvGd3xLGuDXQsxB+IBd6glUlIfZhvO4JlZEPXJiXl5EjLQlojeedySjBuhCnR0cm6uGH
64fz48SUsXlqDrTTW759iceRUSJZAg8I3bGu/VJFM4PA01Y2MWL3cQGsTTEd7+JJ3BIN+o+nIavC
j2YITfgx3Bmmtu5DYpPvyBhbnIwqLirjsGQHe4fUoIgSGt4Qrd7hErngKOemSrmJM96oyPYwo0Oy
gmQc8GmOCPTrk0Nk4Eb/9th6W+xFflUxoyfhhrM2kw+fGIFJpqbyHDWg+CTbLPsDZJ2O/rt4o399
N2XOQPAlMKXMGVrXcVn/8v6yJCvpHcd46uuZ+I7vTgFXRt9C7JBSk4KerLy7zSItxeSotnZqpf0+
8SvQ0wrkT9NrZcChJ8Y/teMB2PII/3dnrguk0F3bTwBm7IUpzvTIyusKh15gpQe1rksbEDT47xjd
wPeIut60L6Khuq3n7giJShFCanqrz2qhr10N8GL6gWWtVXhmabIsSqaow1k7/XbixXu1fETJw3dI
HDkgZASvzBrey3iDSBqLUSemIbEamZDvxbASpY7ePahSS5Xg2wV0QdlaZoE0yuJZImCAD/4qNDyV
EFG2Om9GJndOfjsEJ33hY/z4nvP/2UTKO3CXgDbZB9IGVTRAomIG0h1RI0uJIsi9M7Ds4xujS2eC
GDSqFT8S0BeDLqpw9rHNBOqaca1Bmy7ZZ5vRLvi/J9EQzz0HkWWYdTR/VdcjWNWNBIilV6bVK1o6
4Z6YsPNLzkFTF1AEuymlDHXcVRYHgwLpQ8gtpsjp61p5RAjxqSJ2UbT74y0cb2pe8jia0zolo/cc
Zrl4qCiHGE8wLVGNwPD95k8v0fyKIHpGaVe+8NslpMcAK3U9TbGaDQutPEokOf5pbc9/bamDgSpj
Xgr5wal+sE1rTeEa9UpQbDk47jFY62/AsBh7m+fDqxq8W3kE0ewv+3NyTNFIbjoYRbZw0cG/parR
0UWHZPKvawgCxCFkmQCs8E+Qow52vo/fybMbxJJky8UeVBrOsGXXVza3fy/dsSgRdwzjqWcVkoo2
UV6ScPEz6fwCjKAJB6cNrvpK9K+lOxAyzsVq1kCiygocgo6p9dfI7V3jKQbtljJvJnv3Nwh54WzD
EwGU4OxtLeLCEHREG/+tgvIX6oReM8zTY85cSTKi6nyo7E0j3oucJsGmBZ8MH1Jh5rpHtS0tC/KV
z6ceeVX0wawY47H988AjSuw5HKAZSqH1gf7TXhMtA9VaBBUILhnhR6hOtTpJTlwtonwlPsegHbd7
DOE6TuKvoZY32ZOQo9eL4l8SsCO24265bnsR4Re/zbcL1R2l7IYIotAJAgEh0soCS5/1eMwaX0wV
03xDKatdHxH0RqRW6+5An/z3w4/qLXnTTzXOyIFakmyaC9F+wsYqldRDsxJWEgPcVczXXzE6jOo4
XySmac+G7i52ioLJ1GupH8HvtPCmCbQbdXAv1+7ZUSLqTVdzwh8mzq5xXlh8fxilWcCIdARtZNxl
AEhSM1RYyta5oEQ/sJ/eNhxyMUHBUWgEvkWp6/h4gdmzK/qAAGGKj6lDAbJG8zzdxNIYaN5A7Wrx
Z3/0vaLE4CAKjn7sYr98z/byYzg4HZbdDBZccT3LKC2MZK43Efq4oPWPKqKC0pT6ESGvFDDaVbsT
Xjq/MH1/setCOfETnoisynYQvqlWswOFv66eaTjAOgv2l/beyr6ntrs71hf+RjzbqFtI8u+rGcQD
Zhg75Zq+Y+munlnlbmvqMWTVljjDcev+1h4NYHNjXJ6SJZKhUO6gBXse25NbKJd91bYdh5UZOe8X
SpeLeO9vtqjyRxMkcrqqJce+R/C8I34+8OgChOX/7g4DXCsdAcMd/nsYNs1VGoQ9LPzT9xR1Cp06
W5WRjgcH5OfxA40FBTjNtiTjhq1MMV51xejJSHbuM2fIkUt+VdA8I5etTCszzQpIby0dHgRJmAfx
DjlqYpSyW+ikFNYPfFaO5IK0COn3vZHm9AgjVB7qHjGMKQCj7clVi9pz3mjprG/iG5XsJd8Zn2Pi
WSkekvGXs9tZoHUfhG/zj7aCV2pU3eNgFeSoNra3kxEdGr11CNtEe7C5ROKub0/fstF5QO/ptMor
4Tdovcs+FJ4Ux9+CjVJXBjA6+170gUP0Z8Txk7XQcI+dIlHHOYd95swUQdisniCnFIjdzCfPtWU8
Xkz1oB7CSnluYwFmNjB4sBwQW4Jz/cG6eikfq0OehivXNv2f6mkMGTzhPqHmKv7LsHRt3Hfu19nJ
QAk+QztNYkNspk4hnFLvSJdzwBi3/0G1J9poCYvo8DaP7GVznvbeDOfXKlYoE8RHwrpFHM/flBCq
Iei5Nz8MKRDE+3mlki7Xmwnc7t8o3tKFTZjoD3ztOyBhBmhQH2Zvha2s8Ec3pBmi7T12EDPPjMKd
7Du6oW0TVFl2mAEaMBiw8I+IapJz/kol+eWjr3R+80fok8X26WRRMKXWtILQJRMy/StekBrnRwGo
Kdzv8C2oVHnMbFHlRSORkAo9TnuK7YrQLN/0dYtFve/b0H1uSgH/zLXQqk1l1kVhZCgCQLTJycWo
vwvCL7Xbh3POHE4Spl+ei3BUQxnOtmAeTMnlWSg8wGiJmxkjhFr2qXYUoWlt+DFH+z9Zvu6XQug4
jMQMtjyuBxrt51h4dTQfJD88xQp0UsYUGRU/dTeua9ERujFX9M3dvKeV5LgnYfNGm7HURCCquBRv
EPxkOhZvJTTw1qZ9Px/f5kCXXl5Ra7cyDRMKVuPEdQ+sHzG4kUJ8y4SIAjphcUNCP/iSBv1cfCfJ
G5LPk3labtA1SbzxYMrU48G1zXt5rQc/ibCX9ZTHf7gZExcCIzncXiK3LRZAihIfkFcjzO8fjPo9
Dd5eynzSwN+EWEIqVCHEeWqwXyzLPWsj0Am2iu0xxPFoFHicUaLUKhFmtZPZLL5aW606F1ZOnlQb
9Hif1gj1OwEkkeZVaJJOerualWj58+DNGjFwnUuDaPeq8TYy9EApX3+gytKIBwqGojZtFZIOSoTu
JM5ry1s1pPuSi9a4+oH4QqEg/QDTRReKA2tJFu91MIfOmAjlILXx20K7SZeCXzK4X9JGkoITSLC9
RSmh8YiP7iIz6oUgmYTniOW4r+gBfs3keWUf8A5I21Rn+PuiE7EyU+5ICpr4tlBdmChqPVA83KNu
JmrBw6k93r+M+Cp/DW7KKJZoQ/b9sA0GT1T8Vyf7DDmjDV1A8ToMN0clUS085bRCL+mg1rwBVvtz
+4LeneSPFpYgHaXGOWUtmTxkGCl9PSHESiLgZkaPc300WLB4/UPLfiOCPfGClQutLhhZgb7UWHRy
Yh/RaGLpXgd3OmUcne/pTCNjUFFoGDympS3nu3yD6mwA25KrMJuve52IT5UwXnduG0P0a9MUaJnD
kda7BCZFKeiteXNCc+WxiM1QO/1xT1PbwT8fsBsNuP4sgVtQWYIdqQyiG5dps1GFt4Sm9FCNmW8F
t7IBgEgmeYlfPwP1AxbLn0thips9qk+LCnH6mSbKMaQVbEz778JKDc8R6rPS2olvjIIBxFC2R12f
Op0Qx8ecfp3SGoeNW+4FNXALv+7OtA7LZFQyMhtwVH0//PBpm5dvtVDe4TUqFKPVdoBBtG6BWqeh
Q+T4g5RAhzmHkAzgtDsFFqY0aItZvQdHOUOr31PRd6DKEKTj1d2KJJb1ECGTKQwy8bKSR88l4eMW
/BDjvtcg0nHdwZ+aVYg/GFbJdQWJFmnOsX9TYxDvGQiNdPv2mEUrxE0Vc9/erZsn7TFdxTrN7RPf
+/aPfy22yFklRVU0NP7eoZxc0wA5e1vCFcdJUgYdc/kmur4N/OwVwiSgT5eVSnRMcn6q/9cLaeYB
eypQ+P+xl00QqeB7S6+u0NO6VMPqyq9zh3Y6+qTYeiS5W3C+VfbHtGokZw3/ZGyWty4mxWwI9M75
qzs01Dt0eCGerqOQ3XI/iTHOKrln+Kh4xyaoXtRN68yointoU15WrUnnQ0PTj5hY0Bu6ASxBAEXy
Tdr0lv7supWbykxDBvGl+G/JhjU2czumN6TW1DjkMuL07ItiMIskduXp4Weixe0nqwrKFPGKxvT1
5pOBcMW72pWpTJrdyeB+itz7/TcnKhCkMowiMxB2JuwwFcwF6imN4sry95OWdkxUbpSArwOFmSQL
1F1OwwS5Jmu6sflen2bFf9ix2LY14QjRg6F9R5WfPpYuDJL3v5kp3xUHMlihLYPzW5tTSv7EGk3x
78+mTXxeH0rq7o74sZ7iWgF9zy4qniHGq/jwAI+qIm220Z/jLCJVe3Jfu/+oUEXrM72MhiaCx7xC
YZnimQGNMrfxsBvbDZEQHavZ5QtU2LksrxArOTsDWRAOhZOCHRUpDb26gFEcid/KpL6cro40E2l4
s3xdC4JrPGThP9v05nAdC5Aq+Hi7ZAj671t2qJyxpDMz/+jgb32SgxaqNzghtmEqs79xw9xu0jil
PGdl3Hq9Txdx11wEFDmdUY+YCizIvCNlsH45xHT2Bk9RkHOAoNW3az5LI2aZnf0ezfYYfqUx8JxN
PQNtHh9QoYpj6QwFAu+V6h+BkI1vWFjRGpjMP8qYAqfKC9YhwtAWUXPcAydd3PpvlvUT5WLB/yyR
tN5bHBfiYuzd89QTLg5bXvIPVd0GnUv1j81xB30tYJuotTFHy81RtDqzdcMcUK7dEkXVlwrueIie
RzQ33oYsT8A/i5GAVnjmlzR2u6eCydf/nohyUYfk48A9qGhe515PSXIdRkgvfkE5BgBkPmka7Mpi
PBb7ip4CVCEIyyzQNeevQc/6rEUMF9wpRFkU1j+cW/mu4rZf51GS7d0Bl17anFNKmv222nXh7y7a
JANa33s3mwg6kMUITU1tEr0SKXMxzFiNox8CtEblB022a/u9mzZrDcjECvvrIPJvUfM3NuI2CFKm
4JaiRhX2zNY5mxRM5n/EwDJCP/1uDjV+RDgvg9fTU6ldE7oko2bTGGgulpAN5tdwEpeueAUcNt6H
8U7fRDut53XWFJobk+OmvE6zNKMzWPhO13Xq9JMN0HQJDUucPlnGTWO0bNv3E5WDl5CHmP/wpWzu
OaiHxLQ7b2Xq6+1tNhVd/RsYnz+0Mpi/PUDIxiZcMMY9JY+PGs4/qhKXl2H8RI+6XtVJvEDF+ZD5
dJQ6/JhRSK6NcJrH9FvfcDMyzxqCEEU9wygQAdD6pL+O3GiwS5hBFvq8WL4tHbbjrurnrzGiCaBt
D5sNl8czr7P1Bf4Wed1SJDfJE+sON5Ob7LdCF5wtRI2/KUXNlzvOl832BLeBaUXl8IacSneTQveY
r9ekhZQgv/hClL54KyiRslZGQfJbNUdgD8beDv4Ub0gVz4nsg40q77FM+JFkm7idXBXjqebMCyKJ
VyHDSXqjpmUafxYOQCRGOEo993Cl3IUaEZEzVcMKjoDFD0KSQsuSKJs1Q/H1KUMGfgV1lBZIFHJG
r7gC0yp4BRwAyQA8eenDqovVeAAzPLHfifZbzyOuMLRRHoiqw3WfroyOSXNOkaxYg/5hnKxQdC7i
mXPkok9OEiBRBIDdgNzDLQeSRgIzrx9n0mnbF+e0UtCd3k52LSWDJZcDUfFGL16IG6guBeZ8YkFr
CaWyHLDjx2MNYjLQJxdQ9EBTX5RtXGKeADtkYJnFrcgGMhUqQTxnG1ys8OQ2d+UuUR3cqknsrXUk
Yz6Kj4wZLB7O082TcV24zT4UZmVvGp5cjtDw1HIWQifoinkcQ6sSaG4OoQ9hobClhP1kJa5YNfJr
dUwkk0I8iYRi/zV2eYTsyJW4k8F5c/XnhCyhhbLDosZpZXNVlaboPOkBEefUjyWgyWvL81V0TmYW
RuOSeYT3SOfzkdnKYda5QBKL+HhS5xObHbk3F9MbI17D8oFH3sOwpi6oxQtCl8vps/+3cVyV5e7a
m/SSK3NnZjYVYRosuZXKUu1EeeUrHW3r4ET+0UoXuc8CgwZkXTzqM4Fh+Y7k0x06BqcUYx0TLi9B
kKljYH8KuSPQ0cwEQZHLpCUQFcdc4r1kt/9X5LOhJxdLdB/oJYP2+W4YDoFWHKuEpl1R8LhuqAI1
qW16FJEXzfk4jZaIKRzYo7xw4sySTu8SqMbkczvudPAOUxY9/5sFk/4Iz8baUncr8UbgSl8WonyD
gAn3qbKU38vzeJJ52pI/FbGFnakwDgr/gNuRvD1wZ7omgtEta5hl8b1owObW9dcrH8nAK9qGudg4
RquSw7Z1yAjjglogHSVr5YDGxm78Li01b88bs5ptllArWJcNmnqhRqNwcGZ4p3MFlLS6mu1DRWg2
3tlL9KIG8Z7Q1a81KnOz2cRU+VZriq2P9NHiJvWTH9TtcygPxsYf5hCMDXd49ED/b8W3Z+53ndTY
NGOfAMBvdrl9Nj8jcS79G+1VVzG4zldBMU2NAmZZsdUL8w7mBcE/a8Qub+Y5X8Gc7A0IDyYVvQls
6CWsv/sbGlncPE+hNB3CfN42e8n3FRTsF5eZwojYAB7kj/M5KaBPm/SzA5HMNdKgVQgqGkSLg4Cn
anO5lTbtGpbNPriIsusOAxe9xgwqskfICOCYx5RrncmbQHfxiszxJD37kFAUpd2ZmUJvQv4UV7rc
StniPfXgwcUUB77zsmkpRQWeU702QwUQqspbYNgFOivVpDfV45+YytOUQReqw38wkNa/oDxcOJtx
W/z2JVXTmZwZ3phNe4uoOieGnAmF4+C+Gz3z1twPTmPZlKYFKUL8G9fjC4wE8TT6oXkwyC76K6+1
s6Eh8R6PudvtzUKUQsVMSK+7y4YPkG0WMVuBJAEbH3DZJqRt/22WHohB1oT9IcWiB/tw69b4qcZs
HJ6erro2lLNemV+QvhEB+KUP7ky3yMrd0Y4GyoTe6AUbWqibjFfozTjBusd/1nm46V8TgplM02uQ
A8pGIIJr8jAzuLtAEcE4H7+QAfTd6hFO1beyBAKb7X17IWoZDlVEGpSoOC20bcE2aqhLwsurGaTc
RtNV/l9WgYsz+1Kr4L2ha5PrxTX6u4SJzwgYM3gV0X1GAYlYv8OiuEEQwS4WEXQxcI6h8veyL4vP
Q+rD/2CaD9gewFZcElqRKOXq71zLuMxJ1+FVIqWK4MbFQGSUjHjICmgRq/3VlknxkkOdWRE1Kbok
rv+PDwB44wVvsi8lZRz5Utg7O5aMd4TdEHirKy5cPPZ7h2p+VUo70Zr5ssJCyb8d5/zEv1DARBlf
A+93kYhRN33B+tvOl+zbbqolSR/cEN99pTGUr0TJvt39/TzRNl8tF4PR+FaBG9R8o17u5Xx8yuWC
yw0Y695WwjsmWTXdV9HJt8FxW7NREYyphj9jaz2VJUEDwkeLi2kXKlkkSrsk3p8xY3UsIkgtTW9n
Eu+YVRd8CYeo61TrTrZWlY4pdPdPefCeyp3rC2M4grtqOqIbRkJmOqZOdAirXeX3rICkCcDciCLp
2LPQLGf4XhOTFVe/l+H+d8UHG2xpO3Fw0JcSC8Y1wQ7Fuoy9zEU7Cx5rhTKMw7EXCE3U4j9iyLOp
vOryll770iObPEUb1RcPCG+EZVExOOF3ib+5LogEyxK2r0ZA4qTfHjobw4P8EyzvNE+7ImPIzLDG
n8FN3EvRAG2iem2aRSYb0C+XfOAiZa0s82zwGS5Ee2MKaecIaDz3A+IzjTB38T920di9Z8Qnl7m0
XgXxQoYRKPDBIXtbQmpq1EwI97FRnO2D7c9fAuybuWDl6Tm9G4EjEyj9upTIUSsks/Q/7ZZQRzEQ
Xo8+8HTSax0zN8FflSr1Pivevpec5LNy+eMos5KAk0qjGAeEqGDaQQB6Y7HuLZ2qO1qk4qgvQ/C0
tabG4HApSThOoo33zaT4Yzl32qzMrk7vPjFSGteuWATqkr0oeyNoxfS7G5QSCvXhlP34U6kBExmx
0sHxgxt4usyOsMUnws/Kgb7X9ewJ8ReXSOh5tSTdG/ZgOppjgFZrhWWdpS/9rYTX8j/BXdnVi35j
Gja+I1/fOvPbyObSMNheP3y45jCuXR+zdLPK9ZcIE+9mN649njgwNxhmmNlALa2JhE7qLnczW1B9
beB5phsn1/E9nP8vtJufJw6JARF+spQ1elXvhQnKcqjEasyynzPplYwEhRQv97L1YnXwTB0p3o5/
E53DUtKN9KXidqG8a+433yWvECFBxruu2VlYb2MWs4k5EeKjKqQniDZ3CJ0GLT5D0UGiC/da6O4t
hRLjpW7B4xz8hCT3NnNNZ5sQxFpAkZxJGHJm3CMcXJBcUPGQlVxwyh3sdbKrvEoJKxUoGD7oHbZr
Z3yLafXTwElZiJwzYYZS6BvHXQgMOINst+wGwfKAhypjGHfV4OWubpRlkYoqEVedzdXJOsDgygHU
PPhp/z1Fq4fee/cU1rUND8bzhbS8HpUxAytVx8uG74UL8k6PoPApxngnUNmiRMiA3rF7w5l6ht9m
NvCagfuvj2l+KUugf8Fld/ygN9ofyWE5dFLLzcu25/YjteiA8NL0Zayqsyra7Q3n0YYS5hnJzPjz
bCjAA6LmLMuxrWC4ptG7iyJ/d24CIYpLCNmcDeMQuMtQCjoWo4zJ1JEu8wc8bSTWGkrij5zSTbZm
kmTXwIbLrjSXbKIOAmHyCPjipkKFQavnpZVp+4TOTAlDWyHev9NHFaM6U/nNrMJXiiKrWeJ0x9d0
bHYOt26crznW5OOnNiHreAwpGgVrsglL+TWScEymPP55qf/QQG493qdcodRYMf9GK9CrmxSk0xlE
vJfjvFOrqqI4xGwOVbToIcTj5+iECnf/wzwnb1LU39lXjXgnwAoBKoZeqqzkb8x8iXKKfHdz0kE4
HOivnjcGmjsZOL+zW5ryQApitaK8HBTUSxW88FmzF6mV/d4QT49OvJU5WtpWzSpfNS07fAWaYrve
sTamOM0tDUuJfP9VI0gmHiOr3BR4x1xzK68tGXLxEojV2EHte2GnY5xOsA8dzWtOK9/Yh6Zacs18
bnY+bLpTC6cKoeEoFsdMxbSf+4UCs5L3cpS0NxQo78w90sX/ZEFthxnknVhG+/bzukpUe7Yh6hBG
SE87DeF/AXTS22qAyWVcVzDGeUrg1syB7/Rv/ePDrICxGcrvV1UORIJyx+9Ya+rUVcmx9pQoSbWT
7mMzwYdKtHR1S/+rl4LsSqs7Q6//QtURvVa0hoQ+w1fK3e7Z/Ifey5ijgw0MGIVei+bbJb6u/gPe
2n1nSeSyMGddODOjXeQffYJEQFeJbgzFpC1MlpnN1PwGpGI4p0vrEQbbv0W4/lYlzB3KJdi3DZ5k
VeU+qqD45pNTtLGf2eSf6ZR2YVlCxgPVvOJTiq7+92NB3E4da08GEe2KnZZAcmtidiqzMQDb6ZRn
1Jr94qTWXyf5Z07aU/zpxTnNmPDATEd/bdXHMjqxgkz9b1Xq3NP8bR6fCRtB5fpE/WzCy15gbhQW
TPp18cwMnUlR+UrrAYUJJlHRNO8GDlxrMYcobSymYRELYh1iVaG8jXa9TAXXaBwsJopsWCk8Bswz
24IVU75NCicawXFqBLJaVh5Xl6jwsA3Ezdnf/8zkF1jOqZlesSzKws9ug1nVelvf/1+uCoST5auS
h2K70mRuqHmhda5XI2WM8+UWw6Opuu0aWW35DUCC2rz5yGglElLjVhQ/wJV0Nwt+aJ3rN0kY5kqx
vqEBVtzKHB1uVCLy98j1bue3OZp458pA44GrlA2QuNVjb9GTFk47rYgRK+EJslvJPZoiMZR+kd1N
/Z17BWuUqUVGcy+MY74AGVw+TMklTtG589uogSsrR4AkqWWOiH1/9ba7xJyjtI2O37gWs5EZyTAZ
UhTciFBbzQaKsr47anEKheAHjQ00PW+VBxh2LqMdKRvnfWfZUbpNkUpC+cs2G7zB+lvn4Dpa+HRv
3ZTegGTUqQ+8gqNM6Dpj2uCHq/lCyPnBhz5SL0l2AO+14xyMTNssQP6ObNffTDfAnaG42bmL26AK
z3Dapnqz83NyjeLVypoqPDXpom0JRmPHKXBTr6N+RUdUd4Yz3KI1qpykcMm643WYN+O0W6tBB6cT
sIkcg3N/p+s7R/m8HR2Zf2j07bWpY2MdTeCfUa6p30iGGuAjRjYTM8wBancIgnv5giD1BdAwyF/u
mZmc5Xo2CrKOvAaUEy6Zwa33EahyLgSdqQp63/6IkKMY/b8jy7+UJ0IP2DvGRpEWTbHmQs/i0twF
388Y0IM+oVOqklhEHAIoosnJRtuV/frVXlipNkN1GwFK6kWwgz7k2Mv0mYVYbNBNbc6D3LwE23NE
l9DSblxpLoTKnglJiuRsMw3Tqb2IsrRpvCnq0IGW6YpVEt76VycY7G7cuO+7otkJPP66BAAj3xav
/+xhowVzu5wrvkyCSRYOyd+CIEo6r/YmoS84FNxs0pGVmZgv4o7p3EYmmNFSm571jW4SXT6rzOrq
MJFcHMBKDW/8K07Zs2bc7KsUN4qHD0up4uPmGdhmoRh2385/h1kxagCkqPwG/tMzKv+8/ToxHiJa
HV0hZSmmkkXUhvyB5kcauseKlHeRV3gmHZTES0hYJr0iQ5BgJoHwAGc79Acb4DHhIMhsEHKRTdt4
EoxSG/QNM3VdBipuf4R4c6q/TC9lpSJtwLj8Mp6CwHJ4pK8aqCcLf3R5JrSmqe8/QLqFcqUW+yVW
ru8+J1KvsbbDITTX0J7O5fCOpavIpkMvN7fpKdHmhy9086V3Lnwle/sCQD4Uo6H2rCngg4k6bWa+
60at95FnG8dLrAlqO3khC6uwUqfPF799P5ta0/k9Yb2v0Bw0g2MtRQSBfCNlmNDFhNB7ZKmxuyjt
Fu52SsJM41SDjMnroZ9QM632r2NhuSLUaO40QPXJAYBl5iRvGGb0njWEC0CP36a2L3ZwldAfCh4Y
g084Rolex9QMhfy0WjMtl6NaLGhXWxATqyTUKBilK1Rhy0UWvaTuWcOxMEMT8enTTsN5w1ogKV5K
/WqNlsYg5lhobN4U1Yj3czQEcx75q8UOcD/TzCHM292O0SuvKWcLbvLpj8vu0rzFG3uNTgaKPacY
FYu5K5/afiFltUhHV8ZdgWx1O3CxwpurRWCjyMBxV1PsJDoa5dutm4jXj4LlwXFDwcSHMAqz7I3R
uL+B9EF6OO4byhlCSZY+5XRBMp2Pw7yidnTO7qHkY/H1qlXVe4Io8cR6SomSdJKMzloTdh3W55Tr
pJ3UsWuyiiuF2TGfqwvEXcSXTKfDP0jcAuuVxCvCVFAWyO9foakFhA1TVBWoVycIq2R52EZnu3o+
1QJ+y2HmgGDKTuEVqugkeuY6QUKK1JxIbv6wB81+OYuzSwJfPPIzixk1U90HuT8fTLm3gckBdwmT
O3b71XCe7sAfYAz2B/gHBurutbZrThwCxv/opWIFG5lpSoN754jHxi4BbAP3w98c2xIP5p9g12w8
60EEXvSnkao+ZBhchO0m9QvlpZE8caMlUVYtQaXIJqin1tVb6fbuYaE0AqEukc3+f7n3E5FHbx9A
dCvBC/PM4ONeEGuj0RPDfymjNCW0Uf4ZqPDbLqxWiiB1b0KurPPVcNyFsP3AbhamcvY0djMEP6mU
5dn3sVd5hK2QhR8shT67F8wkjgPhWrZma1haaNKhAaDsrPtrwLWzc9dwwSpKBanx8nFrjmgMrAHj
mbWy+t7XaWrSwY90uoAAREs3zD77X6F7d2q+wzKUv7YoQlwrtu8SzoNvVjQprWlWfbRe3lBrT1Yv
q8vXaOeJevViAgP5CgR+xvkvudS0FAu8HgIcBj/hCgdiCypo5h0QF7u/9xLYL8lFWnK9U6cblE8E
2jIJSmYgWna4vd9yW9GEIUqeRw/zvnn3VqTciCEVAtakPayo1FcJIYY4TvnMu1xiZui0ltTL4RVc
lFHLRibdDHHNzhfiDdCGWSqn02gLXSKWhPrMNvds13HJYB9sEJxelex5KeYATUF0Smk0GKSQsd0w
n/ynMLKz+amawFDj4yhddkoEEFKytA5LDnTy1eyGGQAgxMF6oeCncSHFMxHmMGg/kQgkPejD6Wag
fET181iN50hcnlIUsYhl8ZbU4iw3AfSd8wvsnNlMKd76WA7CQjlQnK9gzqrjBtLSypYJQ9dV3xQP
Jbm8uY5mTagmZ60t01kmsjV1L34aaQ8JjVteDq04HJmIUGEguch9DL+OSKyP0DoUyD9vjQlOIm29
qvwNXs/K8vIch3DOXiejQ19b8/Ol1sZ5WFLR9pIsDyCzQapG2prlcaC68vl2Ckzejgmhmzwr/rXn
X4lAdRR+STuRviFQ6+Br6eXCZ+6S7Q6zU8ElIn/eMGiykJedNK2tcPC72snU0up7A6lAkr6gwEGa
15AO9eWIZLN87wQsb8wkoMpt6/h/8/IPgeXr/AkuNEY/Ry5Sxje4QpE9CaJ68iaMsfLR7TvsCgXq
1iwwseCFVrKSL6qgoaayKQGSaopiN4vev8VkQCvSj9nIMvM1SA/eMTqESfGf1Ip+9nXca99qAToe
qhADKr1Pu0vOPluHH/Y8JtmMwso2WUkRI69wIa/3TEJvsvvTkSppQsbbHb9ijLtqrMhPLJlKHoI9
++iaMF7RhIFUQMTrwvVEfSSnKQQGcH/Fh1P16Qizwr2F2tKOe/5KNbnQ7+BCOHnZRpuC38+HlKlG
a/l6/BZDpoFE9tWUlKWD1GrT4Er7sj+QgOLCOvZp5/FxPHnl+hBKmPeaKVUu+hdwl5tXH0LFPt8k
FnSUVOuLCegERk7tCRCSz5mFZcm7CY9YMIHVfjMKn/5oSOJZmTvGlhXemx1YlYzyvJj5wVbZfHoG
mnoEWnk1GpQg2MjXOJiE6MsCfah4iUyO3meNNd8sxUPxhXpdQTgCtaL1hQ2MSJd+Ie5IeLifHQ2b
hXoUspU21QMCOGln/DpcUWSghHXr0eJNrcHaVf8q+ZvVysM/8ZO20Eqqb2LIWFtyvX7aPzEfsyxB
aTpxw9rNeTEFZJ1oDW4gYGJsRieeCsObzCUTxWPJbUuO5d9sqpuxD+Q9rsq9EPKCjpv0xwKDlW9f
sKwwOhy9tmKsfO8DIWjrRkren+mRaLYFHHO3umOn6/ZAOEl7EbWw6t0u2xEP8oxfDK5emQW7fEUg
Gzrkg8Bp/oAngpAt9WL8xtDrcRIrn178zGXgal+WKdDqWr3TmJ/iywg5ncxHZBljszUJ+lkeZ+AG
UxTC0yGmOZ+nTxJFFkO0Q+0IbIC5zMSHF4c+LofJAo7kjGIjQ+FAaykl1bjnH0eRyeYJGwVlFZLx
pvbv0QpuyXClKde40QyaRuBtcHcxeUfZ/EPGSBW0gMiIgn2GHxrJqlew6wCP0d2O58Yn3fM3xxst
3gk0T2fAfmVn1+NBSdzGNegoBeciK1e4YSHEBhvyhFdCrJUg+bRWhiLZamRXRQj+CtIdH6sy8F6C
k3BYox9TS3lrT54zHTko6xpG2paexJyaZP1Rq5uP0eEYgfz+mkiEI2FDglBG5XtGIkcnr7ayzIwr
uCqFqrYKP5rkVuC39jpc9qAktKrYAD0Q8Ch2DX+pZJ49VB7mgnMn0txsN7KviFLZcBZUvAksHRhc
oJob737q/uTTZwO/Cq+ExbQFZBfX/XzZ22Brv3Wht1MZQvtJdGBRFjvvIFlA388hd/4eN8POdl2D
VDjoW5HTwa3LetQf9diaRbubtghWmk1UIi+priBn3BSxsbV/TWF6E0Zz7F1zsoCT7WbTi5uVNx4e
vbFEt4dg6Z7XBb8GEXejgSfqVOS/T2ckeSsWRvMUCJHsbgIDEovX65EqxtrEFrmwUYO0WAZFWmWS
EOs9DsZoUjDm2RiOEPC7KbTijOjLDaSwJQX9F+wC28QNtUrxvmRJY8M14nQ4OQidGNNCsVuY4cEY
WqahY6ntO3I2kqYVPLba7PDUb2eRI/a5R33bT3tWZd/1xsJaTVhMepvlhOnthig2akz3L5KBVzJ4
rK6HF/16e7xnOBi6ZJbuLgtA90AnzlE2QFIn/AF/3k2GBCX9fxrEOCAY+KpSDsizqjUptaxj07hG
Mnt8iHSQyvpebRLWeHKn76vHb7X4DXHFGjZjtfOajvp7ilkdo65oHD32gbbgTFu98alLILp1OwHa
x1ekuo8MUGEKhXMoadm9w/qaSozfP85drXfL0R9tQRITkOv2dLs8zFzK8NUz7uTWj54OvH2mTggC
uYTpMkqW7lMoJE352ycumPIu048n/reF/0p1CqQZFE054v1Yx6Mq0/ki26scW6S7Tfpl/iZDB0vR
xZ5TEmk7lrZZHWwvNlJCpSqwNEh+5gGJv2qmnUl2rWlGOytwOJJXYsWRkPW2/iy79ke1toVqvLpw
BV9PJYYKi1U8kmTZbtU6XQNWm0ewt0nIMwrJORVLjlHHcnFf42GXdVbzpvvyZ9yqC/5Lq5R9/jmy
3tLXe2Ape2HzfUMtlE5TM3zbyPcBzkPJolOvOR/ngb/cDCm9kC9aX/y0OMBjzKCV+kiNMxFM3VKC
LsKkSM74NUly4+LjxBfMQIyjS6IA/Rbkrw70+pwwe4e5WBKSqjeYIjjwyyzt1mip5SmCw/8W9y2o
wR6Z5Z+i3dF+p+rxEYmthm6ct2ITgnS9B3mc+1c3WyiLD2+MLJV7+OLPNBak22yRJ4LqLyzwwrVQ
bSv96SXHZl3izh6ToPgj0Nk7zie+2+IjFUHfKBfVRstaEdnPnQvpvQ4M30+5LqbzpUvY7SNE3gGy
NxaHQfwGz74i0vykHQIkUZVR7jxHAW3sCnm40h5Y4Jxc/haVt00TSbVawEHtLw3O8ZF12XdIb8PD
EmZfKs/mcPkcNkMVgXvfSFOL+MQ3B5GzMfKAqf7ScevbBt/CGxL9kpnsyRlWDPQpfJin8ZX6dc1l
nKiK/AnuCwygmk760NC3zbb/0q3uOnr4dzicQkBvV+u4zwauxJwIpynif9Z4eHp5DpcqbW7kG8OT
LUxk4Hu+CniRQEnMcvOg49G8OZ5GZ8amt5rWgYlAqpRWQvBYkn8B0RWxxlSz6nhN52adLvpK8zRu
LV9ry8YfxnrGfPCx0QbYWR7dXw7gqLZiw6hL80dHX76yLN9r8zbXZhEE+wvKrZCiEMqgguvNhCAK
R2e9W1Jjm2d9b2wSIYzmwatuCqIUmA2DJ8QNE5TIr6fpdOGIj2mJlh0GO7xzOSFcQk5N/c43g15u
AAqX2pV3YTnyryYZOu0DGjRfJQOF5g9WvJDSyL2MGXSojSnxYSDKfw466cJ9guopmN3EPjEVSp/u
VmmCHLPqD4IyI7v9mImv8z9cI3VMwmdNCSMlklNN8ZIlwgRiUJSQt8MWykIRmXAWcfK9Y8VCo24k
a+PLmytR5DtwIum1G7sv3Rvvyufh8nsSPDWCn1oZ7V5xoxdqWiKHPzysSiqi97iFtjEfuJucWpxQ
B/YMixQQ9Hb2TmYSwwVPwS2chJnqgRWlzlvsSz0Y8kNZYloVQj/QcjvS5LCUo0hHdEO+4n198DsG
JL3NCKA8TtYmOwO2oKXIp0/Tk5G6keqxt9GyUVTL0i8iN41iD1B+UUXvOIwBEDdpZitrQuZ/iACG
O9YZUUzF1m2G9Svu8MZVOBEQmeJQyzVHcmmN54UAdJJ90pWoMIOPPZGq20IRUstRYMDvVcKjI6v7
DSCUJUVtds6fyDhjZV2ylouKOyyPm0nSGhIAhJXtVwbsGghfqr5WF4Fw/zWLDFIiD/LVtea3k4YN
9OKveIMhliB04ot9Y0wfRnS3q4NxSpYbA2niyQ3icVxfB74UbEYe0QCvE8YchEyElYU+o6ys2kkP
HafgAFUcHCUG9des+oxFHrjCRGBeC9w/wMlKlam0B/8cYsckFDJlajSCRCFU7JRcaQKAgK3oWbMq
Dx54iIn7jRB3ryPNn8Qx2nuEkV2G32dNpZqATjJ6cE6p0qRk6ZKA0yRblmD9r9PIJjEkrqe/w1x+
I2WZcIuG+8QGX/rAETsqSQTO1Olg7DGn9AllScuJQ/MB5ubmIAh17mI620EtU/zM5uNocnG2+pPc
A8APp2VE8q3OcUBxRFHRmtMNwUD21LpvBg+n0smkYzIxIa+A60zkfSz08Zrmei/e3Fc+NGqPO5pB
+idXiiGxhCUKfe06BCS4RHZdagAP1HtEOaHQk5xqfzluPVzsJn5uKM0Zulk4Jp8vlnGiDzz/HYmk
AZTB/Gvhdoej655w8tXomIQPutEEb1QZbB4E2fhO3/pfdwwoaNU51wj+5Jm7siiJu80CGFoiEdcq
GhKQHcJZNDE0vQSG4VTeoiIABJeMvHuTMIwpCs3dmqc9WUOBq25nEw8a3c73+vzf8cSgBtRqsgIy
W+Nssu+tBm+kQhCqaKWYA3aJvymAz6wNQb55BauKSCDN64d1hxAkXPd3uCYmnha4oyAHSdaVcX7j
sGv/jhsDM90uDqqJkN26Xyh8rxQkf9+WR3lDuz0Wz+SWaP4TZBq1zXedmbUh/dcgLCTP1nO+FHUK
8OVctF1RHaL+aiUwjoWsUf27NWQ67IjMTJHM9WZB3EaiwaDk8WF5yhjY4LyasFOeH34Mw0rnAhAi
zHsclRuYXf/7Of1znjfCd2OtewLsnUKAJQ77g4PQLNXc57p6d5Fn2TkzhCdn2oEJuV3Q7n4DYChg
mCU2mGgiyOEjNvsUch4Rlq4gdc+sPqPA9pBFYhuYAQCJQardi9QNPH221QKnrLc7NFoZFMYbjsy2
8/Lafpoj64aHpax0AajPQ1KykB03pgwSgPTo6Vr73OoSHU1AWWjrw7T67iLoiEfNmWGa1Tsrq8Au
WEXAxkb9UzI5M45pdcagwarwSFojQgXi9ShV0TAXYahRFgHGvoAA+5fN3WhsWu4jugseH67SG3vj
RLcp1GaPmO5qi7EYrPeVIk6/DJyoPQJDIGnu9p5O2O0v3oNhn+nV/v2hro9xIHGssTdQmiyHNdhb
/keiT/x7EHBUAACZehX0ZP3s/aborkYIGt5+q4fO9AK1zy80lBRrkSSgUZ4R90WBVte30ffNbHfu
QsT3in0VtVmSk/dHtid9XyU6P5R+aBiQT+fu+C7bRTT5yw6vTV3p5ljeVE7AvmSan+oc5q3e/j6O
RMlnTmls5WDYDzheKxTog6ZLSpRxqBTIJNMcDCf0DRklfKl1zJZKVz9wos//Leclmlb/B4fPbrG1
deu0rNzlaD0b3sTy1GH2gOSuyhgWWe3tWJ/JeCSTWvCqlngvy4RSBs7aQW8WS3cF3tSS/cJqCK+s
BCYpGhPHLbkyDegSxUIOIJihiBjeu3ffvOtcYNVOpxi+23d3v5CvEacUmqiWHDLxuX6KsfiFy5dt
pgxK00Bv/wXgSKhvgrGExn61eA4ZEfT9fWx2WeXK31WswVV2mEgO/r4iK7Oz4zRgs2ivw6lXQIs1
BYSui06dfpNI+i7dUFyxjcC39ZYoUUt5HbePAmR/5KgttMbdkT7ZSmWosxB7pT1MoiwUIpgSU2Vb
KT++mV2Mi47UJ85Blh2E79NO6oc42GMuzRvjnkQqsc0BglRFLw2uKkYQhpiFthU2Hvj2lYSAAZey
lWg+Vrwzhk9wBldEdAmjnqegW89se+yWjvC/BtY9Av0vA4YQXa84Vh8RdKnTKP8Ff5jGVJfEjhdy
eOBYPPVhkNJOBrxXvuHw+ydUsASsO9WvIHhgOG+lWzRKMC1mp2twY/atHsWy6/qiwTSdATIVd7nN
8oaLGP12RSQip6DdmgZN1pJ4bY+ceI222U2iiD+gngyU4QKqVMrE/6C5L9Sr+vSljP7rXsHaenxI
hxmQ8hPSzUunpI5EMEmuU6iXIBvKCZOfOt/hGQyAd0sUHJMUWlAKt2ngW0CJNsDeuKW22vnnn0Wx
umQdCV3x6rLt850eJlS4qMCXjhMzTJZUra+y2UnyMR4u0n7mt+cJ1ivGqrGADcRjaRLrVpvKIP6K
n6B3YRBrMSAwFoPgR2PvA25bR1+n/FCR0t9zRmZQ68Pi18psB67BsUkFJfiZwuydmPPYvFbwwKvG
Inr+jsdLnUSPfjQm+c6O381caE+oUpbO9q/pcXt1iiWAxE+aFri0e3dFec897znQWGnOf5MOd7ee
HjYFYC5m6OMkzuPrtRsHLEdhNE8GkgHNnNb2jjbJdCBzjXjsb/eK8t198I+BXsASHzgpMJUDKDai
0BOxWjlXJgG0d41lqlhhjTz5FJkjGHFMg/apDcwrwSV1MV8Ajjtv6KblPbw2oxFtiaJVr19QbGvs
Y5pbEQqVLxVGDwPSnj7Yj+yAm7Xemp307mRW5aJ25jEzqa+q7VW5ey382rqjsm56AnKesnRg+714
gmFto9/noyAZ2u455tb2d6rIa3q8mX7H+ogSpXzv8iM7GWIh6wtv72IDiLkRZ6BM3N8LBOFcAGW2
DGXqmtxSHcHDd/rJLFhzhrDfY2DFm0phZu2O8hawte35TDGn8BFLeEcxs42cyFHIYPhS3MTCYMIa
oW3Weiqv07Gx94rNlpeljycE18/vI37DhYDyYSjNCrP5eEuR8tJpp8RD4euKS2E9n6Dm2FLbEULK
lcg8L0FaZcDM+i4eCfdSYQMTZRT98iMQMw5eL51r6Jv7NQkynuXlszym+RQw1echBYt5TjKfQtEe
9ZtlY75hUt4TqcYUDNaYC3x2pIwecAHf+qgg5ZEPJpzX7V7TWmWtX4Y3liVuiCUIgmVbvSsF/HmA
HAFVre6cHhyPmKCtRJjywA4UOdZDIPr0j2Mbnrody2W6KUsMHCrmQFVApjyqQxc+7wchGZtzssu8
TnukJwGHv7i7owSNQcKk+EOTA0WaRi5OW2O4MdZCkT6EtzijFdwUao1e20A0Q08Zv4ongzuT1X6r
No5wo1F/aQVM+qAlq+hEYn20Z8XeVm4dYPfYmQvkumCyCW+QEpohrtjq9ivD5ZUbTgPID5utg7E4
jYgsWY79sWHsxVngX/SQa5VvceFZqA/O0/K8aTcMCYbSRVdHjLicTg4oRXfhDbOduo9Swg+MJr20
Lv7jg3BtRg4alePhV6XQsVHBxwOxP8jmDXDsy3jm0iIS+MtLSgALEtivThPAJe7kTg+oQ9lKGLOu
uKi+wVtc4EfvU3DwD5KU8mVUTSN2nZKN3pB9QMnv7P4d1oMq1Q2ZCV0g8v5rk5zdeR3jMsuEk5rQ
/x+f6Nxbzy3dzlLo4UzIKEZcDiA/oMt6eK4dKZjv0kGFLQbSgBD4hPqOpGz28emQFNhg8xJ3nae0
+UhqdLlbSO2vgbtB36CtR6K9vz5RweGkvpWoOwBinZaMM7kbRuO1dZqkEPTZZC5fFrEbHHMSJJw0
JbtpvkCqbLOwdXkain2XB5WpQKtuwXNu8T5OxZzjyWT6+IXUCTKjg8jchOrl+O9gj3h0y27SDJ8P
nGLGnp3SCyP7u/Ezpd5K7kLS4qfx/bGRH64px5q8aaX+9J0/hXmiSM467O9SFeLUH4IoiaXIyMMf
Ub+2cNrJJ5VEEuVeOZm85YoMzbae7dAhf8/YBBOoc6GZkQmCKMj781D8TJAm7a/+EiskWyLvHGXZ
i+UP80/O2u5azaisPteimyB3cPAK46DAhV0JZgdVeq9IMrZsDzP7yFiZu/XoQa218Fm0Py8MQ5gZ
iw/2Fbe+AgwafDN3DIzNtHGZSBW3ETCsWol8fFFQ8AbCcHRDQHZ4ZiC/gYBj+Kyi4uT31mOIq+JF
9TVKKC9gsTdP0AVzBJpbau6GzH7PkzSDSXrlbfNkobd6nb2auKMx0OW2qObXIqjjTxUIyq+FD+t3
f6ec/JFyZbCfzdGnv9VVbRspZWA7iFW5INL4K606XddF9wcp3KY08/Yc6bCT5pnuNcUqUzjKwIlB
/AukJap9A+GokvFQ853xYehZzKFnwUS2DjJIAhy5+yDwdKSYVqLXetqSs1n2uQrIYfYB74DzvZ+E
zt/2tBKk7rTlI9l6ZkqwfrI09k5H5MFUQwuX7zoYs/6LNgGUPdwpf6kbMn6GLThX0g8qlZx2ZeGy
cTGdKnboe4G8Q3O0tuORWNmSOJ7FyESBV4VCgYQoajzjWcBfYp5VHz+NJX20x1WyncgEe0Extx+k
LtE12I/mNWgf9rS+aeKGTLxEWrH0yTtpU+Ln6P0jkaxTbY3gF+6toFyqDPY06fBiGTO8EJdy+Xoy
Txg+tBI6LpZgywXWJYOVdDEN6fok7UI3K6UIbaOwcHX+FNUTreHr1J0AYorKcl+anqSvMk39VK1z
vhZqwThN0YlKJTH6ajwvwlheJYw1n1gRz+RpkBsOZIRzXyN0dW0jsEIEh4H/tC5t6y7lKqxVowEf
6Q/Gp5Rr098hn3Xbb5URRG1Idx7ix5r9C0Pa9IjYZX3uI8N6TJ9fccBuqRDeLecyER7kwL6wYh3g
a2hh7pZq66oSbUkjy+QfDPdNBpGqLWzTi7SRqAFcEH27H9MRlCCd+/HZfpYEgIAI9RfdztEQhBb8
bOpiTLYpXWHRQknyE04hiETfqgB526FLBVDHsRdWsGLxBNARo1Flr4oeK1AByzJixlrf+8OspygE
GmW2u5yotmT3nRoKv2l46zM71/fz1oreKZ0PqNbD0Hneu35JiZtI6S0i3pwHOu2Dkn4rS6Qcm3Nw
T8EPeopJ5vb3OTbCL7iyS9Kz0D9kEi69GWXTpQMZn8vcgYXyAOJ00uZULjdb+WcfFaUZePDpF7Zp
+xm51ROOQ0MEVSrMyR+KpZbCJZv3qgcGDUtHV+Vo0Bm03hCCL5HSn8aKLZhc6ItAp/6j6inIACFU
CxOS/3qFF9wPqemSfiX9oPnsF21A0vJtn3/htA8eTHG9dUOPjkXCF2+eJYiAvCdaEyXQw+TRiHNk
MYkd2fYnaCSgx0V1AYa6qm278JgHje18O1vUmdwrB+vCL8Cg5S0qWJFS8xueYiKaPttQYw8aU16u
6B579LgkkHSA3Bu7ZIy89oUpRTORj63I8YC0UV2qczXBn26VfBK6jJxkAcc+uwuU7FuhCgivdLHB
tU19iVPAGkCl/9I/tJuoytifFIKvl+VxwK0IaXuJDF8+P/3rTrF2lH+nteuaBAZJfaCeQVSrv66O
fLAr0DdjB52Sh+U5Q66Ub/b0A+IxUKllZwEiEuss35QAJ3/F5aqhR9ckgn09qax9L/UFDgNQD4Rh
RyTc3NmpZ90bHFlrtMxfEOHWh1PW5zfHgLN8FEo2EjcdcDXQFHWDmRuQ7uNH5iaN+XGYB3N6Ze38
5WWh7XWnxexzVLBUi1oMB8r1qM6pFF5m0uV/YVlwQHTwdZ3orhcfrGk2MBkNa0s+p0FsRI6+WQy0
DvyF9g5yNfH8SBOFZVDWug6hMts8bCCvjwre1QOJQK8ptldfON0qGP/CvdzxN7mF36nJT8135mN3
xdIvJcPiTOz77DLlMN2UzsDIfOEEBSPjKsvfcfvwQkZAk5nRhesCie1aMHZWiL9kgCkkZXp89oc0
e+N8YNgSVUSgsHe7ZiE6EaSJpQSDUoHTLUsEmpAzWkIydVnUIZSx+6mz7OkJyVODn/uSvoVpbkeS
RdOtdEIIE95kmgvjDQxQU2FRNIFOb+JPC6VQ0npB1iROgd5UL3x50EDv5+zp6qRXbvwywnRJOdeq
GfTBXNNd/NeVZ6ihqCKazgN8ZGum2rK+UxT+ddrIR8G4bFAcspF0CPlUu32gGBD11rhAo9gvvpVv
YAwXExlQuoBL2IqYxlVh+QtkHqWM2hhCOY9ApRoLMM1JGgIyT+JD1PqAnthLxugiof6oPMgl3B39
H8ryvVObdP52MtLROjDweGgevetj1Qc3USWEjC1x/g+W0SsZqb5ti/JaSTnzu/yzX7gkUtJkKQyC
+jwLekr3g1WxXQhERBJsNkBEd5l3Ah7RGYtv6igF5X9fXZ+HM89Zrj+f27t9O/glvlbEphbyti+k
0kZiqymMlYKuqACLWxtmhD8IEDen6FTiKk/wIivJhrpyFZ2VQ4wxcxjYjv3OCdvKRt3hwLCiZ4cV
8FOrizaqO3QosjqJV/b0yRi/o5lPYAS0V9Loa4YFS+v8+IDlof26GJL4JmLKGP5KWWS1aRPlXf0r
wZDvxs+A4LC/LuVFdyknQQAMOR4ufNGxg70zJCa8ilbs0SQ0hidBJJs0XkzHoyaEE+0yZkMxit/F
BOwsyiqQlCTKB9fUMYMA2a66/G2D/U/wPuGR0EH7o+8IxinDYqOUnsnK0nQ/V29DUbojSzD4qW9Q
fDpBYOOxOfeIPclGhlVapDxSnwEUkKkIPaNSlebIAGk0Lqhiidzk/z+1wKNZhfXjK+tbpW7rUsiz
vTYKiYIEGqqEbE13UAu2woUyTor6nhWm7PdKFVmy8mfeViK5z7uP+cIiOstJgWyWru0tTuCD0baa
y5+qqElpeLTJVLiYZQYKl0NCJUyKMLF1Tn2I/IZCCS0KPVdKxdnOcYv8isH48vjD/D52ve2TWpfO
I6sVNi+MdsJAGMqqXindvvErWQxvoLgmwVtL0/MgOp2NP/FGNKPBGDg/fmJmBOaUbAizF3THXXbM
dxY+sYgn75yzZT+wKHYOLKGLJQK9KxEq+n4zljQ3Nzke8Xll/tW6FS+JKm4npBEdgvH0f5+KV3yv
MzU5gLuowUTi0TMYhjr7ilOD51tGdtjNsJeLD4YyiEDV4NmNkVuRxmbbrbN2M1iYWtqrWGsLqg7R
OG9NdyajQ8eR1CYZlqN8lKPO1LpdIqxZl3+8hObctwdhU+glsSj/ysswwSZnnB5/Rg0dpxa0fK7k
j404sCOT0s+P8JZqp2eYhOXM5HtRddqg1/aoxCzMkIB2MekUiXFtsXUoMeB43IaO/qnPldtYVb9W
YGH4tYFNHqN1+fkaSGYievHNlC3vO+gSFKCZQkzVOAx3ttlud9grYQRgMnqRJ4mZsZYGyqkYua5x
Md1VV+blW3GBZDgabTLUpKPT7E5+fNr6vFaTXa0QkGG+bM2+UbM9V0kpKpMrfQdNJrVsSgSR4nUt
j8GEEjzoCFNJTpXoLmd/84QTlkPCF3cCsNrt89+Kj1vdcyHtstTFqk3Si0ns6niBK7fd1Ha+0L9l
K501o211MkDUqkVIqYi6KCOG9uPWSvCqiK6wJIFcLH9zMip6cipIl3Xq+vIzXyM3traEGXYN+Wt7
4nWuTxeTnDNR8ZGiS0GdlreujchBuIwWfYIt9LFL6AD+gluhLqS8G1ElrJrEVL4CBqgj6UMS3MFj
C1szaVIyCB/nZCnnzFXWbU7lrgaIWl8PzYmAVMFRTnb9CsJQ/5raqaxJS5+qJ42KWOFWcRPa6naU
HRp+DVbrTs4QcmtojeRBatOAZfDAclodQaYfekNrNSFtT4KkIu25MsP3HWndUpTmR16FgrJ6upll
uqbx1hmDcZdWFiorCvQ2y1y5D3f5YtLk+WhxLi2VvtTE/vroJrIR/7r9wMvKEBc4eEgLceu5b/HL
IfeFleEgZgzkMSvVOSjrR/CJEkZsitvnapJjKlkIRRxTJSZPMieplFIdWFvL5UJWPBN6ZNqQOaL1
bElEo0Vg0fgrWP88MfMBbqeGD/fjJH/dCWaR8SDMgLQog3c4c2+sNqkPbAbIf51EndGfMUrsllRR
AQC3Ea2gJCp1Twkusxx1qDr3iff4IyxyRg42KnpWSTbtDH3Cs+BqFniCX6a/WU6DOPVSxAWD1znt
yi2sYPfVullz7KXWd0F+RLXHujyfXLd2vgmUGavQ/1svLozLH8BSQr4B2ffv51Wry9/QuiG/ZZ+j
ZhA06w1WWIqM+J5hTGO5tBEOnUUiYtP5Huo3joudxEktFL017iZqatK0Sui8lUTfIYf1T+cjPuuy
YBvZ1fmIrNdy57UU6BBWyNBUYoRBLbklsgasfl48nyxJcyQLKFnTA83n6V9XeEMsvUKckr3Pqj7M
AhY0vS//QfY+dckbBTwo0xipAkFERyIgcoQybM6tGsHnHepnH3yMcA6miOGQwQIjCjmUer9FFFUr
DyOOPMCkRmuDXLE58MW5FKhT8K4YWsam6hb921fETm27rhn9Wl4ipSI5zNs5ItEAsqBNFiGyOWAX
Ks81/Rd827ruTApBByNXw5GJJ6lsX4xLD+zkobcFB5rwUQ5JrqYAkIoYAzBB3O5oY00mkie0AEjI
KUaYPR7Fuup8CbHU8OTxB+2blJPnYU0IrKCczqaUvIpsSVe+/qcLC03RD5WP840JBjoPK3YhZYNX
PWoLbQO+vELmxk5rvkVDv7iMwd1C8t6xJ7GTGVYZM38skmWHBraXVuKHVUHMuG5PSZdbyM3DCm+2
ZFGf4M0vZsR3TMiRmM2uPd0M7gk3cYXJ5eSN3naL+tQ3Wh/tyvzR90ZmPFTXSC/uXW3CCBRJ3Qsk
EfNhhCZlozaTRyyL8dzoxhVaYk+pkWzWakqSh16ZOirQJaB67Q/mkbY6Pb7BgGN47gHt/x+eofLv
iaUePRFJfzqVIybMVJ9mSeoADdRpmIp9tqOnXn31gIw2PbL9h67GiJ0euWQnson3e0w3MTsOL0FW
ujxCuufXIKOhV3fYzTg5shtCxfD7pAwYTFRHq0OYyUEWoaylbpGeqki/VY9rkfe1u061U+w0QPVD
P+0ZIhCeQj9bVI5xjrhNe5ekzfxgkvkdlkqOj8R9XAxDxoJMyu3/vqmlfMRFdcnYsTwFAzvRKaU0
LOq+Fm51FPPkWE9hqgyJyNLldJkE5Gkk74F162FZQidiOMzlDNbq3JLwIR5dqq1NhzLs0nr88mnG
HGNb5+4k6vJ99f4EOzilMxSKY+bzEQ11HXDqhz0BotBpNockt/lRrRrYERt68OEYxTldI5NpPtBy
NzvaNyo9rtq2ck4Lbg96hJCsgliUGhmpo9sUTtBez9tlZBvQ4LR3RocGStiL9qroCaw52hSONUcH
HFYgIS+nii3aNsqIa6O/h/gr38kYX8wzIYGLSTgDZrvoPAcE1sriecCBD+7iSbnROePo/2P/8TWD
uH3sBm/LUUKoRlc/IflBkLDFn3MkIB5ndvfRmCO1lkd1OjVd3/oLasqqrCEQKhTN2wGqwV4SBJJW
YpuhEaWfeFX/U942i1p7IsYUHR6sRx391PJHHFR4/vuvwxQRIXAi3nZklATj5cW81Bby9c3lfinJ
LR4Da8DbkUNNGfRBG9kdsS2Sm5L8jCu6baq96XhO7kTLa9ZofjLU6bwK4e3ylwx8miwECO0jwhaz
egOaiPGLssbeJ7UTKNAiHSbr2cDbdHgKt2IBjguDzBlJwbBaKRcr7prtZPRHfgoC343bSn6EZ2Vf
HqqRUD2PYW9/1aBaAea3X9AnZvKF+/vJ10uzeGivLd4CkcC4lGliXxQwXl8ATmtzUEWYtU/Dn4jP
1uMq5dnbCBASFCHEbN6HYQhsymyK3D51WLxZpD+pmYGncpryzgh33AK254qUwiJgbF8+7US0ojo4
LY4jufSmuRjPXGqTdGoiRk6v6prtDtt1xOU68ciyOKVTCPyg6uV8elJTphkyRlJ+5VKP7JuN/WU+
eZlkKztfyCPfAIXA6r/TPF5ydm3UaJrY9Daz6TBPiQ34t9dot0H6gQFIgASEfrppttmwIcCc4q7z
/l2n7cwEFbXhC/BNtz19NH30c1R7zLzZE/5LtXdEe8We/RnsFVJmL0l/XTsD96WxPZ2myvEp9e6h
UdaNiU7Wb0fMJwikh51GRs93g76CS4SHEjkGWTA+1KBQ4/yiFUuJT6lbXtxks8T4N4r0Do0Dp91O
8++C9I70hvjMrT9WzDtBHsh5qgoar0BT2g0pLM7vxH2K1HuRcoA0leGOdWbt4YQMdnynCCdyNzvt
n4B7Hj1HkPaOE3UF4ZarfF2hg0Gxr7tusEgMS18Qjg3j32zBBfup0JL+Lc6Gy37nc5iij9UaKuts
MhoEmL9RN6BrX0sp6nKp6PPaoRGymkb/NlwC0YUMNCCWcQY5WQGZxwq0DisQvA1WRr6d1bIULg5r
ivlo8rnuzmx7gLVfU8lzCyFfC6rIpfA/CqJbaE7UeNShihyoQWSeqpkD+GYTza8oErP3iAQBAtWn
+cdCW8tLxjuZVGYMTDhd9Sa7hXco8MnzvJzZ0XSfQLPj4br0yOi247AR/P4U3tvKHqvxXHnVt+T4
by2H1jZOT+ZcnGsR5yb8qdh+x3kxjTR550nlY7c6RgfUX3f91+Gi6pZtuKGlC2MpsyYzO+A0DN4d
sIx5tFFJyKmEj2qtUwiOf74TFLn5lXS/X+Dlthi4RFPA++cpPjpzdLgckfx/zjS4xG5bWJOTi6Fo
cIBq5uZl6ZMZCnPTAwBLki2Xul0w4WRuROXdgGp+bNDlFG4NQIYP2NZ9v07Vz5MC0MHegIob6Ghj
ffIHi/5ASkrLmUjDtfb7o2ecXSbcBYDmuRSNQP9Abm1/sfZYmRkTtjt89DiWd3ZOfkrUR19c+eq6
c3YhcLrqIw7qZtrIwaWcojXGaxTtsRkIx09ZcQBQWFeU3nrOcebPSu38ehKyQIeMuRtQ1aPn/hcD
VZzd53kHo2o+P+WjP9hapiP7QqH+jNFh9HfJvZJ1pg9e9D7+1QBWdiQfhNJeV8Gjnfff3RH9Gill
I7e4S2BuZyZhvFHwGIuEIGq7VUmmfPwCPouLO2+783Knmi2mVxH8ChOjBRJ+kVDmhyi6EXjcm4Xl
OlwmsVDbMMkvZTN3AHrCyi0/Uwb8zBq3GDXOTc+PnQuPm4MEpKa8/sSECw/zu/zWRGrGZPZWFRYq
ZUt5aJtnPYPc6yJ2q9XNWqzp5C5qtdcWVLOsfcjSCF/oxP3G6N73I0usHDv2w2nqsubuOLyE9HCc
GjTutzJwRTVEba2JjEeNxRyD42H/hJrvH9pYPq3CPoQhr9hnmVqwuDDfSZg+qpy0iCBRX95Dijtn
mxqqNfDR6NXgxDC0/YdFB3FNAC+AUCTByHC/8MDUG/aBkprcx6gJrgwsKE/0qxid4TBhU0K54MKI
sb5zjqFZRXhKvRLeQCYstOtU5narVmPjsu+WNUGv0Gg4tDbooQRmKCs1NFufp+UHjR8PzmrgBXDB
c5bthBYfIOgn8iimi0zEXloqN9OgvHoHmdP8gFHhz8xXZ5jG15pdVj0iDmsZDck+soXqv1XA67qi
/Nk2YYpNytoRxGcYNUKwD7IjHewm3Qwm9Z4O1e7rXOBWSk3CnN9NCr92+tlTdnDTAQA58durC0gk
3FK+memU8yocavZskWM2hCAbz40lT8aJ3pzF9h6CbQRjoQteCqRqT9YcbEFZdK+ZjJm0B6pYsu1d
az27ten+8FbDQt8BTezauwclOwYVc5fMoTQfDhAVVe+JEjbXuoOkIrXjmN1rVoVfLyMBcSUex+3b
MthIFl4YtOhwrhzhCjSvPyfiu0eShmIKmf9IpoBYseUC0AC2oLl12CkIDB9km8T/p3KpOfuTY2wz
fowvSehEBvn5QuVsIdzXhLsvByY5GtP2jN/OqKU78UCAIFS2T+gjQQ3BaqSDNq0p+xZvfRGPN39L
1nKwosFvROZZLGSBoimW4Sd33U9ZMsbKAK1ut1inxgfVeQt7A2uEeQnlmXmI1R/I+DkAyVJJKRJi
zTybCL4OUDbup5jxjcWFmcXf/1fxqx8ra/cKUzzH+CpI0C0C9+r8uQFr2U0FYiJAmXPmohf5U2h8
cinyeAO40AVDwFi2ybzdOIpAyhS2aOpNIGT0K693Ll1VA3fIs3exlHxm1y2KOMExP2Y9cJMhQC+0
D5gkDq+BG7O8IluNift9Uo0plNrAzuAsEoGUXnUJGHH8XIaRSTS2rM/veGdfTEKUPPyW5dfN4v5o
5xt+XteYWbLY5aIWD2xZ6AI/9FkzIX71Fjx1eVkyHUOdSwqlZeRpnwGbdyYm/CPOn1BaqkaKRV5U
IXpkFBhABJ/ttKqk+93aS9bZ6jNByFEvyczGTzOO5X9zqwvUvXMYutdGryaidFut2x9mNuWixRyl
R9RfoNv3OHtwX7ugXrO4wqEBhBvrwe+cb1ARZYbkH+fE8UvofKrPvPwcVW/lDiQm1hV9K6g0Fio5
k+5guGc3KHG0iChnZIW3gpmLVX6XAekdwAPdX3+OctM6vcx88pot/wGiHZ2CpEZuWDhfetJoY3ol
HAIUwI2OXlY4C3JjOjDIfPtXcFgkDwbjWb3awdDxpznm1c/CISdYEtaLMjKo+26d7eHq7voD6UVm
6BJB9c11ElSbxy/PDv8Cu4zttmnUcLl/Rc6tWLSYYoU9YIRj8tsKbJwt74IAXhZD1GdBV+VjZNoZ
4TGrI2R1w0MbMBGDaYeDdIDWQadm443tUVZXV09ughGoodGM/zotnRrcyvkem/R0KfSe/Ot9E/2z
0nnLu9CJTPDpxtk5Wzdf+hHSJN84Ey5P4wPJd76LdpXwKSIXZZs/Kd9vJ/kQBQwDOtNM18iGra+K
0L1MY7sOr4I0FOAdWwdbeAmH4XtZgs3Xh6fUVQ7yKrT/XfROiR2mH4//ftgYP4YWVS1JAKz9d9Fe
muGCoT94OQFlkm9QH4WgHVQf1qwUO1cMIpZkgQYjqqO4jm1NvBO4aSqpeZhHN7oa+hx5n2MXol1W
riqlHnXp/3o6rR3sNfTCRKQrZJo8uZdSq4N99iNVcU/BKfi7iDKurcKJpCBcmOYYfeDDYZECtGfi
Y15sbjIAVwwZcyFQiTym229eIq3MsQagCq5dLcU+hhePPrDJdrMla14ZGiSMgevLsJ0IeMWO5yww
rxN7eXxZ9Rg22qX/DQ1zoySDHpkXWM0L04EQ7knlTF0Iasr9peg0Ia0i4rsg8FS1zPMXIDz5Dife
TtKj861gc3eu5XQoQgtB+Nq+B+iMfHINJegtDXW0NFoavVcvWGn9C4kzak8wpuyJd4XvNw5duNvV
mLlxwJv95P5Nkc7bkWMlJpjF18j7WkFfA+rksJmA8/eCMJpQi045ySbVEQcv065pZt60lY1+dRyA
g18waeZ/QHzRMr5I5lKaTv/ch/OD7tuPbD6ujbDUe2fbkmP+8+uab1yen0fAO1fZXrp5ckU+lpaI
BGAOPhS8hG1C+53fVpSyMn0VGJQt5DZ4zXz6261mZEhiCg5lwK6TeSL0/27U/Dd3aTtLtOFUw8z1
hcgoZxYJPivm1z8d+1D89HWOv+QpSFUUYHBk02u5egP+KcdoNyUA3UkdAq1TCnc8/xJ2V0gn1Jmy
C0ggf2Guattff+Z09YCn6Q1IBKRazwO6fPtXE3Eagd9rFIF6tiUftOlwV6WabHiq5c7ctD7NQg8C
szUAXf+EYxhrT5w0OHsp+Bt0BctelWCGwdnjLeB3+XK37H8HRNAGcuEwSwia5JpbQzdSNu7A/gVv
eES1WyWbqlDvPlibl6Plww6Vz1AKeXMqjbCIG+8bJepnYenlx3eDTNJ3r5TmXERLzzh7tkdocYOg
ZgEiBrkSWG6JhSuZyxvsqHQXnH1eYI6X6FYwpNzLGV79NO/aZQZjJBzPXSAcF+N7G17yPyL30NBX
TOSauu8qUyCGS3FHxvRE/wjyaU3gBxfS1y7KaeyviawQid90tlRA2q+8CWisRjL0/QMN4ptZxiZf
KN0ubRhn1Cs7U099A/yobdGOJY8o5LXLUI37F4gHQWQDmw90lqZGJ3fRo6BeLtNjZDMb++Oar5yh
Yz+r4YK2ntVynQCjtwBzdN259xNnpCstuVjSVKKxb5Ie+PLUsNAqb9BHSbdeovdKdRqv1mLTamn3
6xSHiIxtrjK3+mkX0DxeiuvgvjcddpoIS8KBR2Ii7t1J1HdS6J79mmWR+AQ7gVu0zZQ2Vw8935P8
qQJrO1XHES0ZHvGc1QnX4/EPHlD+XcTHTKttCgZZOrzryA0GquIQRoUMUCQI5iidGowSEcsOe/RD
oqbCe2eomTnpKVkjl9pHjfkU3KTih5N25WzmhWvmfqPtSUTDkWNHNOsG6U2SzvvXtmQw9bzm9b10
RAGx204KHW4WBH6Yjax1RvomXk5R5mO6nbsYeGeT3oGoSTKVyEBtOLCKABG2lCs1zC3hZyXWt5hp
zHhK43BEw1Vke3BRi2XO+X/4JbBVzNibcNiKkEmZausphKCLaIL+w2Uj6ZInuKOfo+CPlkXCxJyG
e3NHeJyD9aZZr7/aWZzdMlI/UvGeUQzgfK/e8m8vuAU3RPll8SlGHTBCRhnX08+V4TJe9SuCxwcH
yYSKOucAa3m5czTnrRo0np+wUmrtBLNLW2m+7yBjdZOttnffz6ikKMgPmoPmw6qTOqlLry/bjlsA
FRkEVxUHAbeNxfwzOnh1dYkAJiSbWXUu9iQTRVSamZsBIlk4huGqAiCrl53DtA8FJGr/UcUPOgN6
r9nsEIC/sOP/zlTOyaH33ReoCujgbs6MOyILA4CsE0ekNfhoUQCRiT3E67OnjwG7hAIsWr7OHMUJ
+nErYJ329BG5px0DkFNxWax5UhfOl54HklRC1W4U9QjhKjAiDgmMrM1mKD3hv4L8xtOFMkHVilX7
EF0E5ZW8QdYh23iJkJhTeCMuL0t69zh3tbjGfjuvfeXnoGc0MfEB88jF3Ou9LY/USc39PK5YBBiE
S1cGWq8UoHzzRpQ3sYLqVPnPzdHDJpyponbV2JZo+vRrmeQrj5bwiZT9cl6syHDH9czbNaMxIxDv
lPy+PYB8xX5YFZDVHeXPKVAUd42yt3KVWWSSZZhZlNOj2b/tHzkaX/HJO7Cko2DUWFCgJfUPVxpQ
MEXoWvR/Z5azsYrNadGnvhgdZ/ffc1mqm0Jg/Z+KGREAbg/L6fVuchz2mn29g68WvWrYVAR4l1px
hRgfCS8B9Y9sI2Q19/dSUdJXMVX3OH0NH0SmDoOFrfOMo80RhYdNoVLo0LvNnedqJ60RibjBLsTY
CVWKtoucXwcbuIHZlwNS/RkS8qEg3OkZ9zGDNdmkRuKmkD1MjrVMfJvgKnhMAKoLEf1SeWI1cobl
lOjnI/czwyLkSZ9BbPv/Iy8VQH99rgW9voA8pf5hss7NV2/69v7//0RKLSAfe6dO3YJaJYfGZpDh
+OaAeArbZEiBKyvZXCSjZHR9ZyNvJeC/I/vDw6XI5PC7rz2iDs5yR/rxv6GiqndKxXiwcfNgCEU2
qTDnpNcskcJSAUruIc6y/s2kdcJ3zId3078zO2gi11ImJ1u39UMr6Ee0QLyikBC0qAMBu6Xzca1J
ZaS8i2CD3y9okfe2tEpzioRyT1sToOfZuPpWoiiQJj9QM6U36n5nXwWSl3vy4FnyE2ZxDD5ypHiZ
XIzmFPM1yik/XAFzm9QR+eHIbZ6kVdV4Myv3mgJj3UaBkOtffulxvsQjx06J2L+ouLJ3B1ProUEt
8aCPiafctPBPdFLV95zf5d3s1zCEE6h/6mxk7D+XQM4PW1zDcq7Qo+8T/beJGl6YADOPcweSkKck
LXSK5C6yB6WNDNnhO4C9bAKmiGP3weeUrBqhQ4joomU/tZTcVzwVmVqFzCOYWHeeyUiCVHwGyt3t
tvtDdC5mRB4TgzJsnQWud7A3EM31mnnwRMUjdQ/J7wEwSPkLV5WFca30junK9VI07xcFc6p5VCqE
tSvgvEsKUZbG6Kbg/+cCIQiFiiNV/15apQNjmrGz1JpU6JBSjurtUQWIf4lgLwurk9X8GVkE0bOX
3ToODKGBz6SgqxQ3Y6syLU83z50SUHfx4QHya4FonewP72cHHFjJ2AFRKQySlY509J9H9/3RlNFx
6OqoxQW+sBxaM3O40Lffqux/lI4r3IKLpixmCLpCtnz+SnnFOpiVoEPmSt+xl1cM73kc0AYPxdAD
YoWzMcEjZwqzzRphsiTKNV5YOU/ZJ8e79tG0NgM0rXRv61i67sLsMxyv0YpvySkgn1A77GjcBx8p
58jsBPuBCWGgbRMm39PEITc+W03BOjl6bKyyc9oTL7WGEbljxgfX6E3GuX2tmPcccxokYk4oQqAo
wFyFHKTD/gNb3fOrIKoabbUuBq7zYc8pryqD3Vr8ZOj+8MMW6yAy+Sv9a1JM9axRX3hgx+bqXw/m
9+eeqIn0HHOgJWp9X5z4zVIGbFfcwEJtvBFAUYrgB5xZP4iIIPKD/iL7Ik7Aqr8TPODcT803OV+C
T/N33J0M9+e1ejbj7MaRrJE8XdPuFzZ+5RaKAVoKn4cgZGdKaNm+CjdNCxNLDup3QHJ+yetWR/S3
rxQ1xQhfMViUNoW1/WsQMWmvFv0Z+R7CzKYyAXRr3JhjpzBQNAygSgtckAQsUytbRFOdZcj0GoXc
zjwb/vmB8BrIV/qh/iJp7R3rT5qb3l4opqOiWMCpmSh9KpgB5lMEJH3GsGMIk7lSvfBZ/J58khjB
h/X04P9Z2oGO5CbPtIWfuS56YRYyJbHdQAWxfbR3znAHB7dU7CfshCvSBg14K3NYvvemIyeoMXQC
ZiiSdnbtGdxOJ7EgAxeAjoHIS6xt4fcK/4q5qZFuPyG19POVtnCDeg5KB+XKr/kGANDcvUl1tcNz
FfpXkF9USssXMsSpqvTtplgRq7wjhoT9CWLo6EebAQHQ78eAwcB4qWVl26owFKsGJAGpfwZ07Yg0
yPRkDb19Pwx+7HvuE7lReMlC06CwOEp0TpJ1Xn/HaWhw9yyzsQkiJrPW/Gcf53aH4lcLKac01805
oAVfcAOiozPj8WYJS52bqskFDVGAfeATo2cWJGKifW3sy1nfXlQ+e/ptW7a6NaQMEbPL1wgANer8
HrpkLZXXWNk5ZwOQ7Nui3kYqNHs/P1aMqJfJddTBVxmr6HLGAAJwubNawq97XTOsU7kodA7URTmq
nRp1jn4h5dNNe2uTFLsX02jN4aCb2yPwob/LIr7GQjyVuJ60SiJwKWGHDrh5MF6Q1h0OstVmz2LL
dJMlB65jMOTn2/BuzdAlzlj+07yz+mkKJzmHucG4LO6XnmENzEc/iW3e5lAjXbYVDNSNGAQ1Wyrt
aPGOT4pujxIzXH6jDN8tsWKvObcR7bftHhmzsX5fvN5GoBv/EFllY9LJ8eVeM531BfvXMT9K8a6d
5/3ajKdnW4vJ2jPqS0KxCUw4RciL9h4s9YQDOZtLJS/gQL50Pv1i4lML/VFCpqoO/hGHCugQKxU+
7IDpKn6Jo0hwu2bU/uwXZiyZsYI4WJGnPIpalblZo3Qeg7MrUyhj/EBSfJDUQscvP7uMlCAIAekP
hX6xGxPcfuuOBbnn3laW26YlliC8tBJ5HpvXXyZXzrKiY08jUKLu3shT1bB7y7tP8Vgl9GAk/qFw
6/JWqovCXIeKfxt8+Zbxf7sRfe7YwcH4coRlgHUEbTKaSh81lrdrns7dZ/pdvFHYl5/+0Yz7G+aC
t1vdquJK4I/XZvibC0eWywgzyNkT7nn7B1HkAN4PA/5uhdTxW3rjCXut/zwkEbnqpfHvEOBJeDKq
Vs3b6T6EeC24JYoxQK+QPrVE4CN340A8QJ9X3SNl9s8EF5jx+6t/8vK3CuEoPSvuH9gc3w9kAs/8
LMKu3OIgnUfYsHE08wIb/kSI6je8j2Blf+/M7XM8sqy7ptUfp9vVK0KVbwVpBu1lhSxJN6BXAKWL
45aFX7+9efMlO/CNjXwrqiliLMaFBQZc5zcUMbu0qe2N8skujsFDAujHtynfok1YCtoaZwRNRIMR
h/FBaqRgo+T1i7Mi/hfdX3nUIWd1kybEd/Oavz+zPKOBlkmoPXU5+7fxtJwLYHakDXqX8/1Usbxp
d8OY6KMyLDK6bBpphMH9P12MtqEHlFwb72Jj8nxDqWGMbgb1WjlQC6BjAlx7WNezPGvcVS8fGjz9
Ac8SkE+E0fe7W+R2d/9O4xpz8KlenUF0Cy8DMvbkZLsg8FfvDtpO9TktZBSjVKNkHpk9Zhn+lml0
7/+FehGRuz589YJX1GX7tJgsCxklfK2DPXueFjSvBvaFT6t/lV5C6gWRAjegVTlYWx7a/KvK9Rol
tZdPvlqz6YwO+VhRuMxhaxTrP92juXHCaLbTyUuXXiUPCc1M27HNRELAfv+ZmuS5hYMc1sdBf1QO
WsT/V3iiUXShNjKQd1gM1lcLFj0OnJ1FyJIBYTnRYnoD+hNmplvxxSBgv7vRO/mdxBs1Xw3QzbFi
Y5wX37OUGT69kCWXbkZz1ZukWFacJ6+W33AHqix2H8SJkAcspCX8iYUuV9u9k0fxtQ5w4Q+F13Eo
ygA+NMkv5No1PxvlyA58xVt0Fx2oYjFvtzpbIuPIPaTIL/XVSbTlvnAijONPC1bFWXcd1CU8U4Jk
McBNdSNhmEfuCbK84QTuq04z4cuTd04JULdyxhGbGdVZAjlz5w1+6Nf2QDtbvtpGhZqlDp0y5bTZ
iD/VdTBcnXwe618lqK91LoqhDyPztvoiINKhs9TzwnnxZe6KANnozKgudXUGDc9agl2KYjsMZyXP
Y9Np5l38KVXjd1WZBxfBVLjJB3LVrIGcEKYGRmXhqktPk/SYwzxPR/b/+cox5IpE8nYVgnpkHBzu
0eR3Z93f1UKxoj0J9OrNiZylQmqcb/mbYXne02kSrDeULkLYSNh5KwR934ppUhzO3fe/s4h7MGFO
gD5SQd14d7JedycRolLEamDS0AadCIsfub0u8GCRbJfUUmRgy7AykPm+OqpE2THewp94sEsPY9DT
x6d2ykQcb9Is20DZyfrXRzYUnMoBESYIkW83iVbGRWoPMmcZvPtueMOFMXZkKA+HJTjharnV78PB
aXcIC3JrakSJ2HiuW2ONoddcg33ifsZ+4DO3QrOqaiNWac/fHsZ34dhCw8463HR8B0Ur2Txb5jXH
+NgWpHUZ+20lZ1g66qNrsnCRM46601n1k/reKXN0JN3eACosbAqVA7vsLxYRcf0JLwmnKOPTbX2I
oawShaPvYVu2xtes14htFSeyDMDrS4sAJ7BY4Um/DBii+TX/z8ovAe73BUoWDqDYxIdTDuI7Af7F
JetNZv/lBE6sOa9e4bu2X3NzeFPVyCxEKsmDHjxxlStZrKxIYdcwOme0bKLa8oed2Atm6/7mXIYx
VrFPo5P2S6w/kfE5TFoEPXxvowq7z9EkBuwgb91Y7CmDnzHEdpWnQNrjEEEn7s7gqU2E6mho/C+5
NWAR60NBXVFN14j/4Q599Aq7FTQVB46RLL2si1h+u70Lw6RRgGBR0AUdtBjI+jGSIzKJpHOh95qJ
rNijtDjr/PKrPfTgqrj2iBT6L9WVa8dhZ9knb0gzPSThJZi0RS+3dBkF3xo0dXfnX+KbzeuTKT16
rUoiHCl6OH2MX4Okzr5GCwBsJZqk1Ms1ndcSHWNaRZ8QIzGZjAblQwk47pcurY71/DzhiLGco8te
Mko1MVCDo34gdmh2bD91lQxFDYD9mbnsM71YoKtxO1i/ihRbaWHFtbP83mQTWufv8plcwjkTpppo
ju4YwTTEWpqvuRakkMP4gKwCIJnaPs2qVtX/df7xjFXpaNHWg3OMElquNW5rpGfNx6muQzbswAmg
8H1EmF2aaN6tv+Rt6nhkmJM5V9oimpyB6DgZ49UQqY7K1LyJXTAL7aR371OMN4KdnfAol438oQVE
T1+HuOKImCO9gt97LXoa4nrP0wgeFwS45FHLVPUtyGm8C0rpDqOWKODaFEmZv/dNuP31A1qw+OQN
n6GFYYSrVyrJ1wZVUHGzNj5rB79yRNhsHUZPPB64GifP7KrTk4N4+0qvsFpJ2ts8++Stp47i3OHu
vhXDPwkOqwcu04da+2mjx41NaW42novvckC43GXkVlYgg1tDy1hnFnYHpmdFDA8y39h5qSq0Xgkz
UALQncDHMXBL77ke9TXhIFKopqsg9XGc6bIOLnOcmK1ofDCl3nbyLmYAHqC4X0JVkPASIv3mm9BS
NQ6LQtYgcEHwNxzd1mpdRvueYYgksX3i4HBAwbSEsIILL2+MLCgpdkixnmyaKzMgcQN6fvq1Gq5I
s433VpnvDv9F68Pj4kdFKYzQdXES4EUeLxD45yhzZCUUt2qpYE3wy4wA2cpc8htVQz4aqZBuJ/aU
t8vvUwlvXRiLHpKcpnrDi2FHLhZ789Cvkj0Peu7SAX5QD7bhMTRixNquGLfKak77Acx1BRsp1yF6
CkKqzsriXoDWfbTYvjPiyXLOWXPYWOjkpLrm6fqqCrVTkwn2Ivul3QO2ZNd4zZpjUSf0SklGdHFl
ZKg8QjLbBKvd9z/ck2R5M1BzACi2ySKVTq/VHc8LvfhltAmxpjHbEpJpP+SnA+m3IFGYqX8ccItx
E9dblKOs2TJyCWC+p0pT+itma115IqEF8tkyYhMa2hne2sQHB6aJA7zzimD08hXys1QfK3IDfVBJ
8qw1/Fvvhb2FRkx8LC1fEfKDhV7zDS3dKx8e9KfdrOrbOaoxshjLWp5I8Rcojj4yvlRnt4E9cj+f
fLlgvH6PO2dNmejtkN9IsGfjJK+xazI2sGaYXViI8RoCpm1ajecKWoy5u6c806gXLwkL4NkM/RI4
FS0zDf3QsyHrhZ+dwRfPHj60Dx9ymJ4VbXgG3VQOJj7dV4L4P30j9riZZ12MOW0PMiOUHvwJuMQ+
BYHsmubjTC3ceUgBKCVUvkVzBwXRvC5eLXEjV+Xr0ur9eMj6ZE7eKlIl9tRWCA2LUYSWMr27xvgz
RqKBbKKVCzgnJdgWJa5WWXpUPenQVZZFH1gItHq/FQ2Ejs1v7UiPWvxm8mCYePZgJ9TwsRFCdEIq
L7ZcW8UEvYI2apwFYgZjGk2H8oQOqciVIcn6z4mNL1iBwZNVEG4Fz7IS87IT0kRTbFYkb+pc4kZg
DYo2Uwm8lAoo3s77tbt3L+Ikd/AJBJKn4DDQo4moLwR9Nup6NTnrD+D0K8Oye0CVCeDdi3yeFw47
riaZKz+QcM1Nth5mxfNDpLPcH+qZLqkkKzmuEUHHk73nKJrqD9kgBie3boRnBkoL2tYaEQ8ZWMVa
lWSMNZrArBpbuSu8ppaMv7mimGHbCaEhA722+8Lb5Utan+DhlOzE3iI/WyfZF4DbX+XW7xraZBEU
jqU9mrqfiJTCwCYBdWrygUMss1qr73ocWv6mpQ3C/DlaHzKLBVEPbPagZatHaLDN06y2TLSeZ8mt
ZQKz3la25Xw6V54ER4X9hIcLSGAYX9lhWn1DvLw5mUxt9OedlQ5Wgdj2diZflsyeBf1rGYvz00O0
WMuNsbnbx1K+zdy1RfFGV7Orb55M54ZS5zFcT290BVQnATOhHvaZFtuyJBO3xDp9AXsdg8D7H1QL
mpcq+gF0MdSYsYLqiCHZMjUN++o6rm3R8i9g+MPxJDwpvkUV3+yygatycVRb4dx/bT+MkwMj8y9B
VBUf1joBgSQNklj3hq7tnItGlzs1Cfikr+6GwLiZ10/6GdLjE7v8yZPAXc9WNdQU7Y8kAGAB4aE9
7LfJt9lBG4yTr9cU+3wm4I35bkOVsRhdMGckDTyshB5h02ShdmxQOzefICT3MkMHSv6mPZ3zqQoV
Mgv/Zuc25Qe7mA3Hzw2sszjZbjb7lcK7kLXulMj12FpiiCQNW21i8P5uVJa/yk2AbCzEHddO1eJl
xwPukyAK2NDMtSgR8m6DncQR3MiNLPOdRQWTTvXbuubUBaoB5KqtUGYy+VJpjWfX7NP38fYQahUO
QG2S0ax/MxMUJTke4WHP8DccPCwYB3N7b3OgRi6BMH1Skel/fOBZzYJMqUGtuwxPLSRC5urVeaHm
ReA8FnkiYVKFCcbiEZbwfTuyuCeRzhEQdvxLzuZNbFW53PEBrEQLwkNGt44NCjSZuavOeUh6ePhM
B9NEReZix630eUZ8Cu4xCej3u0xt0HlxRIFkOi9ZhQEuaNFF2mnZJBpRNHvyOqWE0nN/o0I3UfUv
/UIqEVUFOLOXUZnj0QXteX1amWSO1r6BGPok0T21fTU/NEXe2ynnes7F/S+XLu2fupBSBON/PAA2
8MRbDTz3BmU8NxBa5IqsIX/m6bVK738i6SbTPh3H3Iu1eJAm1fGISfZW+pXW4JHA1BYAddx5mXR/
u7etk5YiBzretcdHqQakU66dOlhVhR0Aycllc2+YECI/uMPJrCSxaiVhSpSn6vXBv/2x2STAXuSk
Z8PSSILduJw9ahU9iNZFZuhMIsZelpdkz4Nxf3TYiY9buyJqL3Dd5Bw+0B5rAfntSXXDy3K78AJM
5+Zpza2dQh7RZAfzVGz/Ssj8f4wukqT+5TuGBmRizz0q/kPCGqB183o9M5XjoTZaKJ73KfHVfTY4
aFkUq/uVxfvQ3+Oj8R0bMnzLx9aZrWPkrGThmdR8Lzi0H2iuMy/8Abx38TBR60Dd8RoajF8P+gvw
WEUQPKvoDscAfYbZ+25ZRAC3XzXvM0XWjZmvvNzFfCGzlKypGS7gyPQL2+vhh9jOcPLHxhwtBPGi
cWyaDmb+Mwvx2/xIcpHDMzFRqA+1BsBLJoirBxEVj0P/gCBr6UbjA6DDqZKHChVCx2b2nTRrBkAi
6jwV8Ln7qzgsKaqjdQ/VTxleCMN/jmYu6u2cjPanUBsMpl92jElGAc1oatMYRnEoDeq3y/pC/09G
2KKmAovIG2fjZwrXVqGbf1VzOCaTyK7OO1phCsbUCicXD4a7yHGdBUcarhEvYwg9zxJ36JIGeqNP
A3YnFjubMny7S3/SnsS4F8b9gsejkOigI3UKqIIDgfDF8AhuhqTvA/aITl7uMLpDyNoEPj++93YG
vz1Jc4j/Vrw1u7K2pK+BWd6laOOkB9JJVrK/UwYP6qCfFOvFCjRjXX951gHlvGb8efKE5Izyybvh
Z7f0YXjOQos0P2XpDC7pBoCGFU8sD3wu5Grlbg4htUouaenFI8+i7Fkyjo8gVkYWTwZBicAmwR7b
5xDrDwWfOQyvb1L40SlH3w+rr3LZg0Hy5wSARTWJ2IMdMldgFqmpegQ/AF2m23Q2enSc34h0SbHQ
U6A3GsXfQY2Tzm0rycuJEbwvzM2lPdkmEklzzH8I8vphxdUd1+f2IHehwAwMmHsaTCD6nalP/TFG
Jj4PNNVvrmD2p/c30hoKeuUdXyBWdEzFncNBjWCcyNGtc0Z/D9hgxDtplqTpkUUJAKYfpcZ3hn+l
QNX/+bUX3QGhdlz3FJrO1r2H7MMase6AtEwgaHv4aQySbJxMl5gOLFj9UdYJAHgRKpY4b488SSNy
0rQjxiifaxKdelfbH8xMxoY/JDVS/a7Ybms7kwwx7Oo94DaHxeODJgtB7D6zOni6cEPYaXvDj4PR
CdeqcdC1SlyvfWlEwxP9jXKA47AKqg0c/RZ4ID4V7JfeeKDLCAnrsLAicP4SpCBhOLcR4178Tgxd
490IkixyocoGMFZnj8HGnXyaQHT7M/vZNqVbbLwTBAmtVUPwzKp130Vc0g8W4/fHWwP+3zG5Vn5N
sw6N0v8NNO77/fRLFBLoYOPPLHNMP3mvbsATOJ6q3SQIcYiq9JYIoeOBboGAdAPxDMtGke+04tO4
I2GH5OkIX/F1QkYZQU6QbYVwSxLo/TJFHOdZTG4+eVz5T0KNYHEdwn0Q/Tib+hWVTrD2q8UfVSwv
nxeR4vrUxSgvwyqVFvZqOD+si+iVuL0SvRAxmZx+coQZkM3rA6uYOthwi15mM/oGYcV8nrtVtB15
nUuuSspW0rvTS4UcfKlf+qT1MXfR3CJImF2eB5ioOiumOeC6+a6HJmPeTm0TRbBUzNkYGke62ere
bIFUzlcXXve4szb9awV3LQ/b6+BBJKl4NDtBNmrTWDdHl92TcNmK592lbAFqjxtjVi4mEiMhIvYN
AU4USdzjQhHp9vGW4WaUYp3bnNGal+pjoMJbu6TZlaVEhNQyEjdDveljlfgG8GA365SYVuOhuz1a
F+qsjsbvcT/zCZMDJI3suVqwqD1fn3XWgl4EhkFbLqHmVfFOSoO5tTrjXLuzMleltWjXpcpg2TRf
UrNhWXU+33TZ83byO0zYLgrYzyQSgrVSoLez9S8o3U8hhRRFFmt8UCVT5w32ULPviRt5vKF0vNpp
etKwVXEbWli2I5s8bWDOOoSWzG8bMf+ep9Z6FvWaWqLdJEyDmuNHr+fSI4goyKrW6T+wk+mODb0H
wiewuzlDfnr3Dgxip2KkBuGkzIafloRaeOnUm202H2rRK0ZEgJA2esAY3crlyhacpq6HfEJATubR
DPYYwna9ZflZcoOki5XJ9XaAeAF+BHXQCV37A7kZ/qKkZ0G3BVOv1OdUrP9xdJqF04zeKa1YkTwz
m1RB82U6ncILM4a8Qxa8LS4Ujhna+FObtABGmNMVo1WjQxibd8fSDQ3CqUUyDLVhlTmb1AiWFnoJ
UGN5uEc8MzHMKzV7p1QgZduqKbp2RBKrMJ3wB6kA6i5vLxo6eXw8Kd+0xO/+t5ClUisqGHzM7XS6
u37Z3jEolhL88+ArVbDFX93oeRkNwEeGVWS10Ws4p9WBWqpbb9ByKocUQcdAIS4c4ENJX3oahjB2
A3GYZ6qThaF55rZ0T4pw1UCxEWB28hocD4qi/fHDmhUx6C85E7nW8i6PRKz44gMv3jVRxekMOt6U
ZWLzuvnmO1AQ2/JEj28Ht5ixiW0DnipaQweqtO+Ei2qNTA1nNvVKKn9SWM+FDv8mgd+H29L8Hhfq
VU+3IPdJTIfo3pDii52YO2Y/c6JKp782W0Uolt5W0fN/Idg+D9GHpHsI3dlgdNTY1ROAYQIuGG7S
lq0jWV+za73KSSf3bMC2ztXZnxL1xMNfUnPzX8bJUXg9bao1+K6V0QZqpx+MLDWyNAsma79a5ioB
7FTsjHMzK1qaxH4FR7S15p57JrlGkGGwpZfsoxAkGp56V5gMsgdH3E1VyFrCIaBUWFaZZzsdzTSI
HLJaYKjx5hrrcc2KSNalrF7uy1aRvohpQfqUEzRKnCe12TfWuSvhTBS95mlwlQk1uDQY2fOas2cd
fW4uD74ZJZgjkMmEe+9DaRPr0PlhMsF9jdt2cVFpU27HJqjGueZPllkvhNYRKGV6eXAzzPwO6tco
lF5xqSv//svs7TZC2rcBFlxTZ4dZvxZTgDYfq5s0CO50Hd6h+AFG1AvhoiQWZyKSCuNfLrse8UoP
M97OGcQDGfgM7MrwaXKbmKpznl7JCrPV3o+9FeX/Vd6MIM068GpQ2N9pqFQJEJr8+/3HLLyaHnej
eav8h2/vmpf76uNVAOZmQCosBgWKfU1/5YnYPreg8ww1Q2GEJmv7ZGpS7A6Qe6Nc/bxGlNSomw69
KBdBhSIYF4HfljgKBknEkcyMAf/E87OMc3+lEkBp63eqAM+CmP5M11QYURhEdi3EQ7NtK3LpyPuc
BsK4jygM0rzFc+zq3yOtGrj3Ye9UpguLLxQfMopZVQV2PGIbTdIySaYJRKRJT3bbWIPfjPzaZCax
8DAyWDkJiBeJ2K0s8sXpeELCv6mJXyKIXbCBnAEhf5FXSA7ENlU0uMow0w+o11gsv+naalSY/0+w
mQGeQCgv2IWwN7f9ORifxr60TupmDhsoDwtE/aYKz4yI3KFMjzsnYVHRu6Q2I7xtog9M/EK81Yk4
XvjZ7qBfMfLpsrLdthWjk22Gzd2W9Jl4XsTN4SZ96IEqE6KjIo37OFR58Y5yVL72L04tXqLlyGVt
LPtxctg8cECuFKlcqW8eKj4xwfcAwFct/xebxl+b4x5QJMiBkpnsXFlHMjWB/p0pWd5G55tmB0qg
gfDUyeKHUF24IS8Z+wYltiMSwG16ug6v7VpUTl8Qo6tM61vht6wrng+MoJ7gcpJp30yHf9kj3FL/
51YOIScmHn8E8/8ZX6opeNXcbVK1e2zJI4IYdpM+ZwY+CyH1z8LRdsWyXMULJOUPLZVlU0GfeUZe
dkvZp3tmGCQelidpUczIQdOBg5gSGhChVbkn7nh9GN8Ip3SCNCnS13k/SDxct2a12JSffmpb1/3/
vsKTsq+RRHA+7+9cliQhxvpJoWNZ12PDTYn9fjzsrVclpu81YWI+cWxuFkySMMMz76qnTtN9q5uV
A2PqDWOqv0eaAuY3qLML9NO3f/gBI2wzbS5hODLSJRSb7JUHdnXmdc5V7ctKEWmWZegMz+OyOLI0
qQpIZAVUe1iCWrlbHCoeY3XYb3j9X8ZS/zAbLhEAesXq8FCb0d6HjBPuQUMYJkWpkNrM3rpy4onP
bU1QJVUsZxM+mPYl2PquSV8+4zbD73aWb9OENvU3AfZt5I1BJb+oodxkF7md1jrXU4Ujd3aN5q6E
+UNww0l6pMfRyXUPaQHB8B4efUv+8tefcByYmoFts/Ix1+gdrHnYMoBz+FDvpOuuvN7kIViiYznt
0kv5U7Zyb0optVOXjnGnJQZsZxHu3sEfXMyyoeVWFbolmclPed69IDBYpDjb4uccCBrbbw9U6VZw
5otdAnU8h2xvKM6RUjUrEEJ/01GAdOQ7gaTGE1gt1GpiSE6WeFRPw37IEGxioC/LStM2aJ7lMOkl
6r9bOP+ce2jYR8i1PujhzECbm/+nxx5+lRwowJ3AsmZ4m63f30JC6z/kw0iU5hNvL9rCWDHHmogb
b2su1CnHiok413yAPh4+CJ7xlJVaUJT+t9t2GzabghevqbmtHaHi4mviLlRJTOarILkUn5Nu3tvC
0QUhebayLe+f7HERlfGpT6UuLVC/uX2Nb/QECVq+9c/3V9O8Cr585F+6d+wxbUblFSa1Qw27HaDf
xkybT4frDJU1G/NlW4JxkIP8MK8VqNzmnZa4qUf4xtTliomIu2z4wLC354uLDrcI07nBweKS/ZC4
XFTPn3P2+9XcdE8+dMlS78SpGffvL7qAEp4NPdFcqg/46pxHalYs3Wr6gfo0VyPIfTAei576pniY
EeYh8gAcoYTeauMx6h8HGgqin6d22jH2HhdQYwu0DtB7Usx1sOv7BEOjBIHYjwBu5D428fIeFla0
ykfXIA2bRSlNEPzI1BZNcUvoNWhEMyE6MBYM5YvaR9KkIiA8/r8EYEKJrEDggXSFY/pudUXjS6+r
JpV5+kd3HoGpIGSKs0pt5PoWRJOUOBsh6PeHG4ci1I9U5+9trbvMecaY5d/qPKdY3EshANjRwuYP
vjWjb81bzfh6zhEO3zaQqctorXiQIPYTN3ElKN7Pakdcmpk1MH1PF8DxUDIXXW4tMvWbv56kVLdI
eMJulEgUJMu6kf+b9lvGs1O/sVtI2cGidD+vQEZFYxMT6QlmKbmtD71ANR1DxQ2bHem4UGtInRbo
PYsBFrqZPjvAp0QFgcA+eoCVH1Ln4P8BA3HBuEUE03xBceCKGfKQt1M/42G/5VmfWZTkDb0iWbWQ
F6jXHzuS/FUGaGf4kFS6MOd5hV6aKrXdIzdsRyMfk2kwkY9O/oooBZdGovn7z0gZs5FSdrXoczFE
9DflTUDC2CSfqB03F+hxo/gcT5gtEHfYF6Ols4wpZ/hu4VXnn/v0Au5unR9+ufeV1ui0lQGCe2uj
zJD/pV7SIXEk1ciscq+SasYosUB6wFWOCj76z5Tcywnsg+j9GRlV0OQ2ienWpnQupTrmZb1EcE/A
IFqqhAUOP5u04hrihfvWFgive8g9G4ocWCSIhiCkpikZyFIItw1su6RB8Z5JHsKMxa/KsT9+H+ah
L6IFG2ExHA2h2sN+GWnbngyAHsRuNsPPvFyR6MG7GtiQS9ksPN23dYcl5fTzWVbgBPXyP3hUiGMV
8sL6xS3YCOk9qfO7JCxwX8bY2o21P5l7E/Ya0mkfo4BdblrQ8kqZ4Ovfe3dQMWVCyjxCYfPqFw2R
Gm8g+80iL/8eQaUrcaQpCF2P0z/V6Q/Ch+2zrhkc3vr7jde3eWM0rXTZks3TjULO7MwowTgydt2r
NfGyHY7dQhveqXnyEn41bcuXUWV3EsE0ymZ8pm6/fOPTg7ei2YQkh4dx2zYKqwCsa7DiowTfDBQb
xTGUs64cCJzEMIfDF5TwPKJjEQZaOAZ5KzRaIf8SsfzOzYbwMsA4x6pk2poTaAD5JktV1aH8D8ZB
jKe/jmD9syfHI+ChDrFiM7ciTsY4ztaYo0L1m4fG5wZeCOwt+yzBV0ukDrUhV3vFqy8jDun8z8M5
rkMu7Oewi0AmqiHbaWEf967Z+EkahAhB1DgIL6g+STn216A+H4/OttjDHBg+s5kqzpFe+zkSQAMj
JhE2OdSQUuadrbalSe5jTE49Pqg5xnZoRbTslmaOAZD9lIrYLC2rTQQj2QVEEh72oxiId0lR+dlg
OTrhNcBb4hk+Z6Vnem3mRUyLwHI64VZyrH5VnBpXyX+cg9a7+yrlXjKGoNRsvS+b/wA8zNc8QWKY
NzLsHL0AnX4mAwerAdSWcaje3W3XCy3yMHG547k00mhn9WQhp5fetAjge9wh6lF+pdUZR2BubVut
Iq2ggmB7QegXLP/oOUziisdH1jbJO0Cbv/8V+xHprwsFVaLnIDGxM1aXS3ijyS+SzUmBcAazkTnT
VdAE0ltNvyMiSpcYLSDYy9OXHtiEvXmem8pgqOTC8DkENwC+49nBFlysXP46uY9ZGj9rBI03qTxc
xzjxAcaCTHOWLA2ElEWBZfU54vm/nuxWmv+cGUPzyaoIibjbbvWS6d7Iwp3tjzkGv3m3/DRIuf1B
Bh7gn1a19q2EdAcNjf7PpMRsqTiNrCMf4nPJ67HnAIPQMQkV9Xx8Y0OhBbcMXbhjKU+eP5qp9fh2
0ACfyLo4XWiQo9qJ5k2Vfu7lCaLHYwPyKvxJKczWCcyCWMueUxqohLdkg6pU2SEVA9Ghk5PqJfNV
xV0LR1/8AFZdiVFe7GR9sPduTIwp2k9CdDbCDDU1zyHtGa3vH+VwXCURUFQZPtFhj/P/sUzJ1iRj
SbEhdzjh0DkE+TurFQJqkCIBuB5mxLyqeKIaC0XMhZfX47TDwJxYXaW0eYWe2Yso79wWSlYWISbF
2SLl7bQlBwz4vNeWXN1XZBSHddYEqA5zZ8ETBKHkbqvo8MqAMJFMIfMvl5Z1HQXjvqPyrylwfAQM
a5Ug8RV0wmT98Ccb4kMsuDXcJ2/uWYOKU2sn4bdiCUqrUgDmyAhYRsRiYycwVvi0fCsEIDjYv6pe
7oqDaHOmDEDaJaPvlxwf4h3rnyroNDbf6fCwXdtvNh7DeILEpKdswo9cbP/bCuX6oTjbvMk3Y4sv
31TmvPfkmUa/3MFr/c5xfsQKY2/tlahVhc66MvHfQfkL2SDcWzqBnU8ZEwuVhWWrs2VPkGSyuFgW
m0V98A8VhYjAihdL43YOb1QZYm4Oi4QI3ULmjyNtEDuMTRDN+334KCstP/AtIZig95ODx6LYg1Yp
ynMeN6a9oCVdBxRrA8wE8r57ppkVBAb3nfy4/t63E94V5ulTpCcOxnAWvTJ/djNcTWuEXMgpE8Fd
yOFpcyIhe3Vg82tLfOYOXhAAL4DJHjSlE9RABFie4atzf8PmZ0Xlo9vbvF6t1iveRmvS5tIAOrn+
mo/nW57HN4SdVgCJNhDaBJZPhtQQj1+MxW6o/6kmSe8//DygnmlnQHwJHkf3YcrRZhCog1qI98SG
095+xyaXi4T69oVW0z2nQcoZFKFxnn8K5ZpPlyYUK8dcXNAYMfhrxD7svRXe4ShYZxhnHdcJhh/u
1hgokSmwzBFJSaUMXq4B24HmHHtXzGgjK8cRZw59Xtt1Uo0Mib5Yu7nPeQ2iltebkbHzS1NtD21M
8yd37ukWapkSu5OpxJvlQo+nGjYJEv2fXJQS0QWtyvNE/MFf7uFg4hzKD46wn+oQULwum2FDEjfo
N+QAVIzPYkYIRBcTesIH9mZxxbU0kP25Wk4uYS71DLW5MWb5Yv71BdtjjauXF4YnhG3M2otNsy3G
FsOC9qugLwqd2pVfSo6j8Fa/DdL3LbHtaGJdBr4CnhdA4RkTHgkkFqWpOpg6gA0+gkDsa0US0rQH
53Gsj2tWJX02Ry/uWMe/SopD8dfNJJxoDXRNwgAkrtIRTn0UYLpNlwFhqTYm21jXzyu2A9OZy807
K5NXG6MJHE7U7mqQzYlTjiO+1//6chWQmXpId3ODWKtTgsduTlMsyu1Nr7FroUhBr61rKqvbu2pN
e7AH85fvybOpyzT8NwDtHshOTcf/B0u+PcBzoWv2YZzsStj6u6GBmbr4o7YCaQSUA8z7SrkBqEHV
mSr+c5RcWNf1kEN+a4VyAzYRHjcJZXAFKKXyoNAptyNToUMZPm//gUJ1AzEGrmzOiyMMwNSZnb3B
l2ZzRPEuDwdRcqlv9+fM34TZ35Zpk+mmVo+rKYXl438dH7Go0jp9AKW/1LajI6pqFQASJO6dXvqy
TTingvAGUM6rmfXLOOKu8h6Uc6LrLZ07TmWsn4qK/Wdi9+RSEUr3s4HovEQWBELQX+tnsq7OfQW8
KdsFYfZ2WIo48CY3mrbsO9j6ea6vMJobmnUl3XLpdi14AJu3bXAbO7E11+tUPzi22DxPASqZgqXX
TPvBG1Aed/wwC8/nd2d9KUys9ORw4lR2JD/yRFabjcDtS0lzYPtM+HyA7gbMuKRncm7ghNUz5KiJ
aBD0Hxl0hlssApXmMG8Lu55lP+h2Rvge0+vGcrjTAy3DzvXAtYVtSumvNuyl/zLlQk9pbNxWEdxo
E9hmel/UPYb+5NVsTmmCrrw5mxDM3DrqtDi5tyrkNZWjB4Bx5J60qDUoqlNTNyUpjiJKpTJZQ0nG
Z7iz8+pz5JRj5NOfJ+Pc9qxwZ5GLgbT4w9Q8GMo3ukFaaQx8sK6rFlaveVwTLyndvWtxsy+is3mV
14PSPivWh836XgiaOSVn53hElx7WDFD7Uw3WdVwpyZyQV6+Jg/52JKMxFcOXKGkmI+gHXVkR5fki
bz2FFg8PnDEA9o6ObA/RfeK/4Wc1N3V881T23foY5bURKhRhh8pyg10pbTGtDYkGj1Cc16uL3IPS
EZBA47Elj7CraMi4SJx8Y1N3iQldmajzzfRdiLvi4KqGROiOHUvwKXKU3IqyHlmfctYCpcurw+Ba
D6jhmkYIYGFYC9waqyzRnf67Lf4ym65gAAaN5Eg6U+W7fFI5HnaNQPJ8NB9FhBi+kQzhkAd0RH0M
XbQSEbafRW4eSXd/aQQDjGe/B9k6VPbRGkPJRWqt24fjbKJa2L+WGw+1sPeKOoCG9L484k1MqaQY
VSI/D8ih2FuMVHs+DaJCyviR1QN8pfCbb4m00OPPrnwWL/9S/u2Z84gEjusFfGXhbYb8QJacnUCB
/AAX+zNJKVxAgJFgCrKKGdItHxbZg1KWal7FSSO8Y5In6k4lmDiXNyhNBkwCY2h/SiWXjoPK+X3h
mxwY+VjYy9PxVSQaQPYUezbYpPnQlUq+gmI7nT+gIkeHI3SrPZ+WGURdlgajGQRal7lzpTvjZw/c
pH/PZeZf0YCu9UwCsq8ZbtIbDqmf13avVVHmsHmNxlHjyndpL7Dy0+xdx4WwTbWIodZxUTp2Hmcj
edA7v6YfeNLix+bkymvOoJkK/qKBui8I6ACndnCUcWHiyMfdhZPlnKaFXVyN8nluIOLl0PO3nfYe
gTjz77RjuSP5nGv08Fni5d+6kaFEQE4ppq16XZDnCqt3xnvE7s2DDro9EL7geURoQ/CrBg3TApsp
k3ehLqDzVvtTPZJJA2493zEG/6ZGJ2euMHA2jxdLnIG/Q4knsnNIs3bisbCh8Vu1ivLxDIfbO2z1
adDIOkhvizwX/jJgwQC2sJGWtnPMR2+gr7S8x+NsK5w+Ut9FfheKJY95LK6FdyI2dEho8Um20mHj
X46DKHqXiBU9IMmbDlO+c2j3xJX2ULq4PhIA7OgbNl+F3YW8oLTkWQQaako5WYw1DAuEjnHapxCx
4pFuAELEHnVJ/pXAQTlNsR8GnH72J5Ad6tTjW43g7Jfy6OawVTETzJYYA903ULZbnG7J/gtONNIg
yfCnxg18LFOBHZwioUl56zsrbPw0fNw41MnpCVI2kIPxS2+sd3m67GlaaZCl8Z2vMXE7eX7LuAwB
B0gQ2D2vHZ8sQTx3n+C3qbF7Q7QRiLTEFG4xy8eg2no7ddH45zTmsSN5CAvrYD0BrpVOcSrRXK+E
r52phRC7yG/RimQLse6ple6E88j1mM1JjEC9/Rw4L2xyfwBTPnkl++iZY+eEI2OJ0ag/lG9ItR8b
VS+i147Lgx8HCjgXzeYYQdAa6dRrWjF77hQAPzgyAs+sN0eQ/12LNZzyoFwucHgGwZqIDkAH+xbC
r4r3N2GRBMGTl667/9853+kKkE5ouB0hTIqDAVZFUJA426VaiUMmNaxntUXHZA1ZXf1y6s7fuhxF
DjFVjOChWqqtwIyqEO5CT4OFzUrjhtRY2yKDHs0wWya+GhDCQYVQnkFrw4xzf25ct2zbSWhDb/Ji
bQIqMl8K6GzpmEQLy98lN1/MC4NM1c7sTA75mQfdOGyK/9zxINLY5lfpuM+SafO+q+323rQf8/no
voHr476PJiqB0UqCwizmDwBS2p5r9D2mFqoPeQNGp2hhYx2bTYSdrxNzGR1rQDrKbWkw22rY0qwz
zWz9RSZHrtATvaib/Iy2qtPmhGUjdtFYA36ow9xf3a0ACKBh3OTbyiBLT5GGbYmOU6zopWy7ouNs
xJ7ewUKHqMjQ3dVvLDR0vYOS7Ywi1jmDM6vxLxAyL4Nf1KuLsCXFn13pguGnJh+rD2JD+aHuuBvL
EGe7v360y/mq4RnG8nuhwOJrHYU38G0DBtTlP2zbogELJj6y8NHkrHP8VxnpeeX69AmvUG7fnbl4
GJzNmEkMOR6TiTZyZyavBQxgIUHRM5HX5VklemiimxsQPQ4kCVvehRfEPnQkpDNkyCndrUUqyQkx
ePyVYbLOkR4tn594GxHI6YdsVmMjWk+as/u4DE+naK7EkAGcw7H8aDaMxs2EuWDZ7RFxGftPD6kM
UqnXXMZ238U70Y93Sm2aFj+UGH/yJkMyiJXfu/jDlZKecBdwJxIYrF9cvZGOgihINEMWCXc+M48E
+XGoEmBerxIiSgvaEr2mzAVmW1pg73AgLrHozf5ZCoGkU2seE/UR5Ic0ZTXgp4JCWJWe+KzlrZYK
g+l7n/9WFvLmAfYPjEC+mC+oywF9j2NWFB6MEdhfdMf4wYxEvRPXTXnFX89ZiMdN98dCXEwQmnxh
uZf0Pcr41p+y5JAGZPS4Yda6c7uanc9Kc1fx/46cywVMiNKFPbuNxr50RHbjhoXdIfU1LLCXtAK8
MAWGV/GgRCvl0ujaZHuJsnFbA0henSWJTA2grYKInkr8/X+TCVNMGTy6AnQfrMjYqyRRVUztnWaE
V8QdOZDdMHOqrEPpN3CDRF6YQ9XYRSSufLNgJ+E9neEkaUCp3+i4kFo7aA04n9StAe4/v8NVMeqW
xgqBfPGo0z0piS29H4NWap9l5VEKQVk7/tlgr8/VimxjzaHW5A5Ndyqefkv2PtU298RBEeS0R7SZ
0fGUi9A/Z6on3KJVLh79sVJ5McSUUdl5wHpcfA7yxcW65zpzmDx+21muToWEiP0pG+OTWLYxDF4C
nRlHz4Ya/9a80TmOKJYcvfYgb8AytRMIeqDgm6FbS8k2rkKj1PrODnvCA9xOQ/wHkuSevtfHqFRC
FrvNYDprYcdCJQ6eu/76xHtPZYe+Gcqy4ESnyd2RkBLwtoj7fW+TyAHOs8wtd6J2n7JPf4jfeoao
cnt0kMmLeTw03GHfCeqA1i8SqK5EuM0w3YaV0jbaUMQCaOiwnQ3dK4cea8iueeo2o9gxyVchb72I
TORpf7H29GBnURQuwufMVctlzHYsDrksAaSMxXpgglVIrkYRXRrOXTFHSUZl/mDpL/VySD3Xgdw+
YKqE0I1VjkWvkooSXFYqw9IUwYsduTPJOIeJRyXHzdaC8zAjwaSg7gOlkV4cZRGH907tGK6Y2t08
rUzSl4o765kTEgLtD/hx6/e8hLIm228f1Vb5CJsI2ci/3HmyvE1II7AcxVfndbUzPkVAH9KIwiDl
h+kcdvwoOu/InaHyI0v0KVbQWE8VcJeAK4EGz/sFNMuRKao+pAx6PP8i0UYlD9AgUIolD8AuJVpC
31G3ugtKklCTNZvYdu2zvfoNsVMentq6kNWw3lSp/wcId0gjkVPRgjBFXmh8QFingSlIoj6eVPYO
i7BkvdEnKSyEA1J8m8NbnlPVGD3rZruIOcNY8EnCN6sZUoQFJveWe0mrt3s7DPrAfkitSjgwz7PQ
1e9AtgQRRZyhNP0+kR5YfrZnKpLQZ9Bx27MgTtem5eWJINGrXsFH1lQ7xUnRpwRsKruI1TDVL7cw
MIyWPE6ts5nTBLajmPEBV1IcWBfeaMj7tAD/PN2msEBRRyGEi1xuDI5pDpo9B/ix6vwBJczuuykD
RzghpO/n+IWlFBfav6Lotf6grP0sq0vIH6hiw7MJa0bvPEtY+iGfU6xQAl3VO/WOOq276nUSJ7ms
2/B6jrjcj+SWng/p5YToJsVjwH5SAok++PewgaNIZHamIFaEmBB0uYQiOWkRiEhBsJnlP4fyjxmw
uqN+7qPag31xd7wb5AtJT7iUbS22i4KDv/rOd9fdpReK1Oxd3XX0VCI5gtKTsy0k9TrTupO0F0Eo
+0uaSdFo7mqaqg0s6JMV/5NzkujFR+swin7Rzy+RiLDT4+7Fj9LU9oHKipsZFEWtKtqvITz5k9iM
08Qu5nvynJp/mEJRG1rlKydXPOk4E3xv5R4+QC009EUw7kxpIY+xCHQAp/uXWRTVMgqEq6Azjhoq
SOyHZW+FPFjnDjJVhXUkItRv/MC27v4tHxq83vgTP46hG/63q6eizPxrooj5nfGN9q5SEFKvBGCV
wa5QvcnDkLHWFNl8vIoPQ3ehc8Cw24bWhI+wta58lT2Q+wwcQSA8SkJC5eGzCMV3q+y2TOqWJOLN
0NqZBK7WpDS+0ileBQaVvGWwH0PlYR+ObBTEJ0bY0k0puR7LdkW2ZEcbcSTdmGsGWhnLmiZXIce/
maR7Oe3wJhv+6Zw68vdCjQr12HsuJ22sgTchYGGZQnhAC9VOUTo/9yV3X8bBF8o0pGbmhD8YBwt8
BWf+c2JpT2NnWYPjS65aUHy7bg7FzwBwQ730U+u3vNvZNFLrEQzwobEu3fmlxb99phMeZUWgAO9N
cAM+1BqIfmqzcYNYy4TriR+rnDh7wJ8ByG9j1v2h1Rn1ciG6aKP7PVY/mQ2viVMVGV+dJ6u0BSm3
wV9iYBSDtXIFVPKpsxtyTPq8ekn+/FYVX102732w/ADhTPBWdgmgk4/3CVkHrKPFEBkPfPBFEk1d
Ge7hm4/WkujqUhphsifVonP9CbF0PWu8gzbahzJdkfZBnHoEAEokbyH2Ustvx57H5KhHz59spzN4
dY1zb89BowclzCms+QvFuFrLdE3xPEPYiRYOWvD4LOl28e/i/2cTiHCU83B5P+dWzqn+pAx/Adx8
uHBUi0awpa8zVNQuqCrgzC7+555E6s5RcEwJ/4NpcnxIN7CGNKxJmQx6azFbY7KdjrwwFvlMsHLh
kONoFCJEw0oDF2Ir4AA3vwuKOwEKIQi21RQ66kd1hGE674BmrxgZWg/Eeosfi57kbxcq2o+I+qZh
8R6/ku9jHgriqU3nc67wm8BFt2bcjvcrMaukIlc/4d3pIZaHS2JuwfJ+tCNX0SWq6lCG923JdmOS
CNljhaLkizBiOphnMNyHo/SL7dGXJc2OBZz4xX/ENmJxIEAIH5I6Bkg+TavGWPhO2v0QBCMk3UUL
7VpHz7V1XOjYjYBCBWu2ueA3Cvz/Zbd1Txa5SNF6DfYXXvsfkBQ+3Q72u7u+VyaVBxim4/Xj7ds9
CYPpRXWk2Cub1/PVkyaIBPehmxt+LDnfTxbLLTDSQpfNkGXErBE0aMI5mXVagNWxc8ORqg/nKf2t
6VnnDFU8G6yzHweNAPIFgbn0cFwU5p49Uxzsl1V4yMxdu0M/JY7yY6MSFhLTgEWGhLj22/jVRYXt
cnjewrqaUVj9F2+9GLLdEzmfJbhWyIWkQKYYjl9P2ijKpzHVVhzvvAzhicjwBCZ3JQJvzuvYsvr4
z0hAyYfpF7kLMtGhcRh4rNLNLkUhZ3cArdZ+zug/3qgQzmcdaXf3oGzEAvLRX2bv6OALnmZBaHaf
nXtVCXp1iAuB4K/X4tcd6uCv8qd9mYpHu329b2Lh8upnDqFUb0pNWSoYE4YwXpwG9fJEf4OJu3Su
+ZXlqgIeETYCsumnz8txNbOYlQMlXt49ViLpy/yyFd1FmREwKM64xJdpYu2r/DO4WQHgFyH3m9Vy
93Gx1ixVwcAFKo5rDIOrQ02VTNSZ/TEXbi5sgdPLcB4RuXCGcIbMtQEVGp0fF7lB6JMwL/sjRiWo
N4Ix3tIsEBMYmnD4w7zbZhfw2JkaAFNEBy3gxr6KPaEikUtAP3dBCNxktlRLjdWgo4+qeNRRSt/R
/73ljRc0MNy1KYPq3+qT4V30ZLG3951GRkXLqA9xgAeNJkBanPsvtX9aTLXgsCdgyK6BBSrKxV6j
PO2GRT8zDgqnfZlRG/v68Z6ovk6pdPrFXFeq9XktPKofht3mxlIqp9U3SXNeaw5iHLzB835E1IMM
vywg2uiDg9Z5SXchSv/kdm/0L218XKzCOI9Dh0lgd5y71qPZ0NENlnmJTtfyW4oSNy8/dKhOLnT3
JWqAFnjXu748o99l2WRI534IxcJcrAI2EZxTxqc6wHXIgyA4eZlmUdEMe7gq4vgN95k+CbewsRjH
fWNwDdbUQO6sdnoxrmND6p3aj55HXWq+o49xVr4LIjdLvIQChkwYfIy9bWnzNTFzFK4gM/lRg63l
lbBclQFR+mKKqnCFnwf9cSTVcdaZQmkEsHmb+9/3Uf17mmSUgkRS+HAeQitHzwcB7JqbVyyxp4/z
r798JO31E5Rl+CexFCSa1bMriSIj0JOFzG2zZoOPIYVZ2KsOaLwyYfRKvev9jqq5RtwsSsgGElZK
Xy7CkK0cqJeU0aAuprjBolxeK2j18yQI7eaB3o3BneXDBdq0s7s0eoHpepdEGdFBV6jJ3g5iTXwS
QMqF+Dihl+zAha3+9DQK2gEkLYJe39PGEJVYnTgikjPuozzWGnUWP8UdSg+JBmTqXMYbx3FcfWFs
i82IRvGxwRw/lrBczK4xQjp4RKRfnDKzH3MLCJQmEptGw24+whHfnnglXWOYwDwAdgtFMj7j95fy
zBD9kb62zaLY9dkMVhh7MgBIweu1U/DuW/6Pt9BTMKCtDBqx7cN6y2/W3fOch8uD15yyOXGfz7k7
t6q8aqCbAGUcNr0tE8hnRZLAhH/Q5hojDMzTswzQR3vpAqEP5Q/7i7XpjPCfQfWVkCg6YP1vKFTA
Upy/wEOm5TmTPERAY5jtk1YI2wVGpzrbKDGwa16gmy0+MMfrVDGZEbQhLI5bhAsJ2uVjH/MDtaPJ
iXPv5IoQm95FIJVJNnTJPURdeGE2HFaP7EHy9BE+XzIv1aCHrxKKjRZr7aOP+6Xlkx5sAn0IH2+u
3m+yaxJzjSaCov7YJz4OMYGdLvb8UpAw0mmHcXD8jIEjSKPZI9eoUft8g1VpXehSUYxEidjLOjcr
3enhu2ML2pd68hvmY0TNVZ1dodGwo9L0LEaFuERmTYuDXN67lgZqjjh1MxzBNorZi8XLkcTgVKkR
Q46/h2/12zWn23lqxrt/GoBqAa+vpkgcLPNyIBt8sBBySKUDKNSoTxgWEvSOGMSWijfZzncJJfMy
YWjV+fxfgb7OGbzQnKIJVMGMTKGT55itKdMYo8LwamiUGYMIptLc/UCW8yoZfK8SLGDT3PTZ0b/a
u62K/U11T795XOqQx4VNwS/u6Rb8sLYV8BMIwaNhe+yJwb37J4gYxu++9TFZLABhqYrgENoyB5g0
q9knnw8l7bB/mECXG1EoJkeHdcUkCOzLPrULZubmEO0/+Py9qJyGaXygnd41CAGjRHXpIPAQTzx7
65urXpgwTe9GdGGXPBFBJtfyf4nZyBoRIkoe8oH8z/AM73tiZqt/QSJLPJ8XVc4xuOIlvxyCh8aQ
CWH3d3yQRiIdqDvX+SduQ6m8tK8bMb0z43U/PYfXA/DTPIzXIVvf4pePW/qBdf9Jtj8cCQiBYexI
o9P5yK4lt4DIdR9Py764Tt8k+KJbADL9fk28y/Pvt2mGrysmecqAf2XgUAKhkNM1HikpgxBnOMlJ
0cA5SpKqlI539Z91wMokYr3XxLGPIdPvE9XxSxwFA6Whvtv0cPiJwpcJfI3zfAu/4YYBS9zPssp6
ZNf2Fr9yl4diBwTmavks5tSax2JWx/5E+HT97g6Bc7iLK0LZyAZiKMGEB7nzfv6VObvSQProWtW5
jYThClHppveGRPWIAHixLbc/tFANbyubq8qC8TCMrpp942YzeW/unhv4+EgzSvzRqJx/W9BDQkqr
XFo/Bjf2wt9HzY6sv2DdGPpTdbHAJRcaK5CT59fTQefvQW/H+G/wiZU0nUxnjq3WtXcOuTvk38EE
pKO61F3tK5JQDAV/GwDby5AU47fX5VcoBQhozY7OuJkkoe6//xWlVJjkmrPaFSBIVVyDlwaZhkvU
arQR6TuGP9eohQdp1og56oEvHAtiWNV/BbkdFEy1uvAoixFf07IrL4lm0g77sjnwfuT2LuQpT4+A
Dzmda6RcBOSAsvFo4GFinoRq52n3qNrOE/psKLXpBQvv80dy3JrUmZ9GmVG4Tvh8Cn5DULzLwDIu
O6R0GMUZv9d7YwRQPnN25wzcVU7dXxMe9mBKvWdQn+fEs1VemjHbBlfIUuSdhKMJyv274BiiR9fG
hKqxRpXDmYeBlO4oDTfbqxLycT3NG35ChiOVQfwqPMfe7Lw3umL6H9uv5/I5jilf7CRCY/W3cwcV
1o6FhxKdz1fgRmsq29xp+mt+Yw6MhK1fKGNe2rbft0JBEakiqaPUWd8XKcTxPEVpq+geGspmu1Dg
Jme/lx8p1DWI6yTg7bMpz4A2C3T3hzo0Tglm8OqxSCGCwn5T+yZX4tmYhxfxXIxK1d1U0grhHJoY
TQ/pqlE15rHuCqH3b8uHNnYf2mTiCc7gvH03SQsScv8YBIIaamEYStIIkfNuAr3d+jFfb0HeuDsP
G0egQiYLVBXOAncSr5ybfCNfDjG1+bD/fEur1U4J6TipZFYQ5hZnoiJo3cvry+CkcoGCvcDMFU1S
+e+Tj+296s1j7GljfWEQurRDPEL0rSjMGHRbhGGiDFJSa4GVuLBzJe6oYZSOD+4/xo/xfJp84Wb7
lk/+p8DUfRRJUUz9bnlue/Wdj6HVYWpsab4hz5Vm5oVWlyTZgBRlUQotzkvZjZPHk95aBf9X4wUh
UcwkK5blr4gYVH5SiLiwzoreJn0OaS2voXpSUoA8MkoxmfpzwdNky72i7AqZ1QBtnYnNZnRTsEw0
jQGBk8eo1JRfjB+QDERO/XbuuEjYb4IMZVK3ZmJSTcAfXauhb+BJKnmeOY5cUnYkIPdBVZe/A+Aq
fhbF/NBHAcp6ms35QNwcp8FgeEWaUInfPMmDOIND843u1doqVyENRuG1D4LC6xyuC5+qH917Hr+P
a0D+dJ4rsciL94NyMbVyKlddKbWejelpef7cNstAm63ZB2la+/iuyFyQykD1BIgu40WbDWPEXJPQ
PPuoEFWGpdFBCxwFxeIWlj2zbzxjV0ZFkcFhVJthgX7UhP98dwqCqT4naPACFidnuSMuZRU4T8Q1
+98heZkaQDB4h2Ol6TZG+1YMkTafNLZvZZugZPhPo+3XZP864rsSnMLfjdr+AZblSaFad5v9SQjG
AnyvOjGnC1el+u0ZEECDv5fpOPIJBQCiy7FDoaNW4C66J0wH9vq3NhDqwGmXnDTyaGU5dv8WyXqc
EFmY5bMPICmAZRRW7fg7PfeXbSVMyLQtoxECtp4mZhM8eURK4ZlwsiBnLniYxd2Sev9PBzGWQ/vO
0T0LaAsxMkUerAlpax1TUYN9JwUcLhmwZO0rmLQzO+M54Uuvx/yG5BqkQYXQLiK9bEdNPKo/yE+L
5spO3rAz0u92lOPrBYJRT/usnUnFhFE31xqys9Sz2Qkjwc2mdf5eevGWBmV0KAdbwXXuIwTTa18B
UWoHnqQ8hVHh5ArFzJXTMMdz4l1z73xtvrrqp9v1iKoNbx/lxW/1OqmIdURiIntM2K6zOJXdZTyK
eI9wvmeYyp3IibP9ccck8DlPpb4wi5T3P+ZnyCg2OmHlphO/9btIRHBCtc/FMaW9iYiyk7BaHmP2
cQB0g9ngjgDMLIH5sOoa8AjSZr8OPrnk2UrObg6B+Sst1zVoR29Gs5QxwEyzC2zDSbrPLxf6VZZS
R8J1WNQuNNG2Nl+lihqmtZJitWo0GylXpgl9DFTw6X7XINUCVj3qgLi/cJxXY2p+DIIyi2J2Qn6M
XH4NG8ZC6NTaBwyF7EdgUC5ThA6wfoOGCT/kPb4UO5zK+jZmX8MTIZRCjzebGuV2ZsMJ+8DHyWHJ
COjSzg/3gga+xkimzhuPby7Q3Lzvx0Q8CvxA+TxoJwYN3mgmpq/69X+ahJy7IRYaQb1ZwgOsMTJF
r5rVx4OjgMVJHFJcfDqKt7IFT1c1XPBrk8DFXl9lqQQBPezzbAnMMvIbrhfhs9/vS06ENJO7PzNl
M/zRccfb3Xy64EmMqqwiAaqo00m8ZYxg05wawZOJpIxAfMy5lxt7+27Q9IlH1dpMWwPL3VNqHNOJ
ZvNBC9LR2ruY2xO7x35CJzEmw1Ipso3on51XEEu5JiVPrhKEYsZc66Zg7rZV4xbjF48Qmud9Tz9S
xAH3VtPDeUjnGQ5RoDVLBZzToYLgWlTPGAL8TLLSBQzlJXCC2smN050ZO3fh7vCVlNeqVsC4N3QH
BYH9BY3JtL/DN8vXCERJISgJEvyoAAI5188sNHnvJadRvq2V6BHmARD9J+aDPaVGsofgvWw8zcR3
aGiyz5dJQWYtplXmCijQ4WqCUa3a8iU3F5+shtK4jPdMbopHpBZtBeHi8Nfs5J7EGOr+b8r9rZL6
oVnOjzFSH5+U4bJ/vHSEYoWlV0fJFvdAeb6diXG55EblYRiC82hn1mXXE2lVdsRSMRDprfseocG1
PtR7m7zzVdC2yTRgGBRTPaEBr7ExwJUSZRiHEBq0Txd03PuQ4J+OvCABWzSvk5Cwjld12sSRl4xB
h0d2g47Oy4wqAoXhNOKYPLgk7lzeeOXMvRHT1I5jd/sESMsVMNVxi/1nmRfVR5V+X0f//w3x2KEA
4hghv/PxJzsCNNQW8zocUXgOQXkt5gO8wELfgx6X5RhzZKOtvX9uexMOlmPJC/Jyc0fzOPBwCNSK
iKnAAUEJM+hKBt7ICbl/juFGGMXOx5PdtXGsy5SJDeAUArUUUvgZUkspGclSQifHXbdgBNrGQ5Cq
KofQ6K9OId6MQOocS+j/2RdT6iDYj4Aor1jX2OHsqrK1E+yDOCgjYXj7x5iwUsgpQlf9JPPwfKXf
WNql/EdQNY02t13poNCUXutvlYLxxJ/nxu1KLP6yD2VAiZ+GK4nYyog543Jvl3sU1giNPNcT47ri
TLAaFg2pc6s1nZeuK/552qTQqhHMUCaRyyc7XtWBcocqdsuFm29s2hEBzX/HP3Z3LU7UzMk0F2Db
TAE5o5LeLd+HhSu9/0IfMAp6JN2pL4htzEtFXQAg2513QmIYWlanENSabZBNPgRRlXVcRpYGhM1l
6YAgeRGGfGZfgGl3zwbYFyUmy3HA0xh57tJTnaobQyCRwWUBgHQQHBgBhvuN5YK3ytd2U9Rgnuro
OPfIBzLfLIQpZg0blqNP5SLv+ggNsM/YCiwvrcwh7VE2bTmBiYGKj/omYUxcshYSzrCzl/RCxjzl
8LP1uTRsqJnHD0l7Eks8aTcGENDzHQ8NQdPMEL7+jKqjsrD77bsSuwYFT2UbCeOW3ollawsY9j9v
6WmkugxABZPRkyc/b+u+nuoanoxd4sdqY8+++BTP2FR7GJgqcM6Jkf42S+drFH0tZhAtklcm08GC
e0mW/o4UWGTLi5OFqApqOVPqAS0307sa7SdNQ4ERx46HAzFg007hRRGAJlfZQzKxKVpXoAQyIZpk
rm4hwYMXOUHSk0ZpZkmRD2cxQjyjiUVjItlcoUJSYtoUUpYcdlP1BDK/FlEimyWYJ3hikMMMIaHi
ONJTHKKDyPdcvg84OD28VKFIuyh9QNJyvoY8ABh2cY6OUH7y9FXWSvHwqJ2ZWIbRQRCQjUOq6fGz
v2aIVi4p3DnBq9x6u72DYkVv4BhJCISE/VBaduztE2eZYzzCh+bUmIwi3uGT3tBobst6ClWP063U
vkvpkMDh8MQKwZYKIgCrgE5m0TkILbscvfGJVbjWYPK7LXYltGRl+t5cUxfQMgvvJq4kDo9y15cm
0i66T2g7555EVRglhHH2wjY1MszMBl2EZI8omM8ovTwsuS3Q+9FStGEGah5NOHeWLbn7ZEgpsOD6
UxfGkTNsPl5x9FsIsd8kT2X1zdRDJ15Xs4KSmMLIIGuoXf2vuE6A2AajhJA2CEs7IYh9vcmSnXeu
8rQRTsQu1qNorsmTzig21gk+TJjqQrFfwP6bFMGxfLLAaYcbi5OiJo1Sb97Y/aTQVzumDvhsn/Z0
u0uN3AwgxEVCdd1kpBh3WEG3vf2Ke8bIlzZvcYjUHG7L7Yk0I++hiqxslUZ5o3qdTsTJ63+zuv3n
IJGLrJpRHRxsSRMxuOyINptWdIPu/rLAMlurgPMspSVft/hzNzI6dpmvf8besNcJMD/Lq96U0nOE
UqsXMmiqcMxJqlir4dL1EdBjMkOqUyEsAIhMQ6qoGGhIhSI80WKwKdOLSaH/1CbsTron4gF5sl+s
omysU9mOY9qAfKyh0AL6o5aWe1kaC+Gyclpzd0nfL1D6QQqvc4DqAZqZbM45Nv7FPkU7EGunQ7L1
i3oGG4n3vsg2efxHrYBPTqpQTCK1BuFgGIusuJRgEto6m4k6NY1cFwqbdm8WUam+tm3cIGM09RaS
Yb8VKM3yMgcewnps2R0jnzJJ57tGu6DBCGHjV1fLlnVpC+O/F4OylW49pz0a4z5gTb+W2A7KoHBA
E9yGOdGfgH0LYAzMCJ13jUnZAe0ILkig3K8Y0q6LrWb0X8HfUyd992bY5EVsXz+wzowPr3VW+h8q
Vy1Mcl5ZG+Nq0Js5i4lnXoLdDUjlgueEW4Eo3lN1H/fjgKzIdg5VagpXv+c3FXKE1UTrE1cxFCsM
mhqWxELwMK0YJALef9iT2hZq5W1L7kD1pe1niFaDMin1eg3CjvD5pE3ATJDyy7P//i8PDlGZi//J
+O+cc1aSqFbilC+luMW0PGwaS2+vwzi+hI3oo9XcRoU1OVFtyulf6QFFi7jucW/g37EHyVwSO2kq
bKRmwpFQuZcWV6J5T6Z549npEv1BWJc3qGlkBdRaqwRZO1ie2cmL1aJ6oP7H2Hn0pg9ya/14+10t
setYJaNZIz0dJTyUEGUKO97gAofzzKeIRKbAKHwW06UOWx9dsZ3KWhucdAW9nD8A833QtpMYtKh9
gQ19Rpv/S0azwh7U/3VFgCi6fmRyxnyc3okcemoc3FHuN1HR1jbzjW/IwOl57vpME2rvy+EQuWLb
rVopIw6jPgZeMWmqPdaGf9SrJDybvssJj0C89qe/e5g25qRqG3rWmlTHIMPsjWCsczznT+FYtEEw
G/j25PGD77hUo0nXZnhJ0rO67l+MOBq7jpji61x27mmAW8iLa9RujjYYJuvAAKoCyVB0CWMF/clY
sKPpBdXAEVAVZpgdKUXtvu1DHRmKzMaQpTl+aMTNcql698ucfXbkn8qXX26sOEa34ZsVOiDwFJHN
QejtEl2ZRnAhObEYzY4Gdou2nHZp5TQpG20yjeNzL/f74VCVStSKRgbsdT99e0dbwKquUrFmN2rS
OUbH+lzpRYks+LIHnawp3DzTBNloF1XzL6Q7I+dvXJEnLdX2W4VWR4L3PPR1or4+2KRXwKUcdaCB
nfN1Hssbyfs6eUsAogH73Uwzeodq2abAP4SOo+T9nJHd4bTPNctr/EVaibQo8T+0jNclZQU/0E4+
sygITpoXGtNic3gOAIwx7ZIyuMV2mbH3qJlIBtJn1NlH7weEXOhs2RBu0CYerlvadb0Vf+iON7MU
ouIBhE3mvGyjxcLgrDwf6WxA2EQHF/9pfIVHSOdSOcOE8Tsk2XdgsSaMMh3OfjfsTnkyeVtHJ4v3
QtFGb01lUm5aJ8brYCjTLfB8YoaBdIfKQ/HbFjHKKEjHzZf4QnE3Ytx2uw5L4H5LyA49AMUOY6md
OCRO7BzCihHg13YbBc92gzFGMPt63/5g3P95TlEbeJWhl4uljYtvwEXTRL4ilhnRw6lJ8ZlOPfrP
JGeTK1FvJOE03aMa/WH/zIbfOHh7v3m0vcW+P6SwFn8hdZtCMcdBdTb0CoxtyMDUMEkl1Av5rhgU
QvC5sCIYeI5MIGZNp2mYTFgV+ygPcg4CJ5lAa62mK41xcMBJzVmm22G/8WAwzkP+2YairXB+1xTg
fzibd3hENFw8z+dc2wfsBsG6KNMcGXUVjv7h6RC6pzw2CrJ9Llnt6VwwIZenckYy6DVDxuQ4+myD
WWwkuKBcUAfL9tg1YWk65VxagugUAPbVoagAPO6oEGvqyKby+ENeCtvQhNDwZwht7ouKpHxHchx3
OYGl/F0vXS02A1H42Yj9yOCYFXoFFSOHsHQRL2Uk8vTYnFc3QAnv+QEMfI2QLQJcO5QqmURvLI13
7LjkGQOn3/wHCUy0UjbUkRws/D3Wi7EGs5ZRzuUEnpNrCxXqjzLNUPVfHiRzpBK3t2lt4c8kG1xG
XBIbpAyi8C2ysVUJE7Sw0/9c3tvuC25NecnFVCxCB/e6fKUu0K6ukaCVSI/L5OVAxGrTKAAAZfm6
FfgDLZDwXOv2IzMMT5iZ44X92Vh4uL8EZwr4Q7Zv400q1/z2dmtplco+4ckiuDBYdqr4gsvJFQWR
JeQI/3tg3Vz78h33RAcHZRzLEx50g5IPw2nbgGOw+H6UOXvzNu7EhSr92Ql38wrrcljTcD9+Ts8t
MSd0MdsmD8EFYs3JevtZTc9tBsmETjpgqvG8X1Ny+PP3QmATEbBb20f+pqU3SgwQAkYryK6L9BQi
v4E7MQuBqSOOJqC3R179JLS7QMHBaKAKg92Y4vfj8JXc74dj2S78mduMt8Xj5qH3R/q7rJ4bzHnV
9suqfEAnE8QiMMkoGTNfRpALBliMXPmhN7H83krBqCs9Z49V8wUfBRbwhW7xpNqkXIMhcwYnloCn
qx7Q/X02PP28WNsi0zRVErSMbDkwjAtBhAhB6XFtl1aSJVtddzgD/uIpwflVsPs+6Ob/Ydr13R5C
mvwltS++pYMJzrnTsFJCUj69ktlWR0oh3HxdPZZQ3wCP68ex0ySWLpUQn9/CMmqvsT0nQRk9w5vm
coQatv4vbIM7sIJVMO2bk2ZC8jnhdM/IJ7ZbKM56bP1a/6DI2YgVkI0tqzYR4jm98f1FbAcBw82P
JUqX9aT51aGhK04WkKevEVPiGA27AWZl5VHL3js6sOSTJN5B+8nmBRSytMHmflTaCkcATu8OLY/m
5K0YKJTTZQQjAjsXvdtVfcBPEf3e3oUNcA7pDLurab7MDvKZIYfYLoE+7A54eFe/qx4xDW9IR8HX
6G+wtGH3VNl92vFqZnoTD6/263H/NdOziS+Yysj17POZQs+LgtQi/xW0OD01+hgnN104nA26cBhm
SH0rmCTtalumRIlURhLYUfdlklzyvI9VQ1i5NBWONlrXi8DhKY8l8EEJKyO2yh6yux7ixROD1noY
mmBkm9hkSt82jYAm6G7Owgpxm6YWl2lk5ic22JfVtOnaweC9VEz+v1sq9cT7y4YHRYZfTTi+R77d
rmFWsPcKWDDkn+7BWa2DynND9W7y784M9Sgta7cQdxrmi8rvELSmkxP4Q3OKe8OWhaHdOUY+jaKM
jMO7R/GTnHeLcPeF5arBhT+ZtR48Jj+5e8qGCdUg584dv2Zzf1ZEe0/BApD4MFVVOdpwY1ccEt3/
R9lp2pzfHKI+V8ImKVaXtYF/VWLRvrje2T1p4RkQFfmOC077yepziB7C8CgoZt37eINQiPrSyJ8X
U2i3J39MgdDCzvI1iXWBoFQjzu7XMEi2R3rX1KIWVMreJRSmPD0LwQT1fnUK1MoVoFcELgv5AEkH
TgYFLQ/dALmd2jJJDZDyasjbNgxyf0chAYO9cAybn5xrSSIISjJf5OSp8ZQQ/A7Wpyi89VPZ5vVg
kpiQUbSwCO20EAHLKYld0kXtpKkkjYGRN+MfDu5JtF6UyYA10KJDGaM5L02E0nd/XkEmbwb6ktcL
l9OC8J2g9VS8gHLHr1RaZvhXzCmaL+hV+c8JmTQ2JdeEv2Edgss+urRDg9+uganTjPcxB73CX6NJ
OmaEfsE9aTwmz9kAcANR3ckn3SX69LJim4R7yecqV/eMkOYvgmPYE9CfMqV1LQW92AqMbap5gP6V
vDQ2yGGbIxqhpn4pIvprq8tXMX0UufBvM1kPZeXs42Ula3wGa31kcs9WcQSENgPLJvk+zBzzu9Rr
vPNh7tuYVO5dZn1Bl7PilM+N3Kx9EP/jNztKbD5d8A2M/b4Yot9+r7YCWdnhCA5reaa/kzcVD8B9
Ju8UCTsfSxkfemWzb/LxTGx4i9W7uucF73cI591nzpf6oTWSC+VBbtYIZu9y0tU+I8IyD+7MAyEE
QYVmMYhBLESs8VSJf7ZxxsKiU7C1m555E04CnLCKXA1F421LkNWSRvfs9YQvT6ShByHGNEHt8Q+b
ilv2Gv71/Py4DxZdtuhA/J0uIsQzBZuf+7Rbh/ENWnl5ug8pdp/Ysl8rXnxVE+L+ACT6TAJFx7Fc
OV8V2ZdAryWKP/pgeXqYULJRox9zN+ibcFtQzFdw+m8/IDmHP4HoNJ371ucxIDGqfnPyHE+1jjKM
PocOpDsAUxHoYlqjN+cu/zPYvUdswyi5vAYDpDEfjP3tBMQgV26hQUYOmPqfXO3EDemZ+D1dk32r
N3aaUxFMqg/Pw9BHf8lqQWdysOB/eZl5KxM63EAAmPeXx4kmRFj1RRd3RiRjnekJTFkyvF2DRXGS
8xpZ3nsY9Edl3AxJ3bJqtiSnXFYdJwjmjI2rOFMRftL1M6PXgon42TQkGYRkHjpdp/GAO2cpSYFw
QAx1CDw9TX8bCoWMfHCro3FYsN0DBzONVlMmVy0svK3NaxgLkcPYQwSAvQIYa7GzsTJ6CGaLtcSD
GStAxtJr5xlSCLcDg0AUv1ARlK2Dw/I5cZ4jIC/1vekR5M1lJfRmQi73DQ3tBlk6/De+mOU/zX5Z
5+30CsDszQh3EhPWDLPMnEWv0YGk+GXH5X88FnLVGKPuFmAU2QtQlOCcG8yBbJLHlPazb6htxsMh
dIWEpUJo5VEVC5gkFsQfyMYpMv75UaI8wvTt1SV381Q2Cegr4VCBg0O99NV4VKOxwCIlLIPGZBeI
h//vGyi8fN3MkeJuzYyHf7/tX4JtyHYTf3nLv2kvr1fr4AH37zlEkMVnigv83T1LU/K2o+kRqCG4
kRsDLY4LpcAFZBe4Y9HHSbY9EaG2P5J4ZDpA2gRxauO7Rvkm/OhUVGfGk7RPAX2Z2d7BITrh6RFb
Enu7Usk/QbbFbLYhr2Vw06PfoQzkZzzQVWL9AV+op98GQdhsCCfd+JRM9FezaBR5xjPWQnW69Hkh
5GPG6XYJloMxZ4QfH/oT1qmV5kDZ/ajQ5T+qKu/222/vCwp1wHCX6uQqilOEZCQiMemkZm7kbwtd
Tvnh/AtaujR1etkpoKmblSAXlUjyUSPac9Pu6DL1iVwkyf0uLrusfSLGa0nLAnZA58j9O9bkejjn
XtIMezRl0AJyMRfrnyGH1MK0vy8gvIwcUhiWaBJJsSBCU/T/oa3G2FBdmXAhsMmoYRBgRW5U+A2G
FHB/G3f/SDQJmkribhcLydYQH9pJTXMicwnAKThVkZCydmiA7KztbnASrhns4zRGRo+QvDmAIZGH
jA5eI25Z3wfRJLUQd2Iq94aEs+V4z6rEUlfc2fjlBFNiGI6rx3663azOufZfnF8bQmM4NlgRKGuC
Vy8/uG6ZEi05wzHCFvfMPcumqV46QyckQidYdCr1EgxUwOT+3ZwvQzABwh7tJi5n0SU6Sa/tlm6e
dv4ffhdGZcdFSGo++WEj1bvIz1xNAilNOgOmK6bVSHi389RuaDwqQBoNtTEcwx4Rn/L1k5kU8Xyl
V6IcFMY/UgaugIqFcVM4QnCz67VOSKQc2GGY5UvBf00qkNjNoEMh5ehSjPTkc7gx77lDTsVOkipE
wNaBRNpyWZ9tE1kUmCUIDrGk1HC8FChG+DVDgbuABk7AeXBlATVRsxYnqyu9FGFe3QzGcjDb9gps
YDj4xZJzD6Mx20fbU9PVqyDCWk+8SH8VevUp8pnLWR8ICCcmpfZuIu4iehB3Y7LpjO+QhTX1jLtw
61V3azNfruw5W14ADOzxfTbvTJLAfT++l3ADbiI3u1zQwcw1fhb80wxOEtu7UHa3REzbzzgSF+i2
vi11nEm9YeTHsn3Y29Kym63Niysd6x9Drydw5y4nvddLm2EOuhQKGAyRdWE/SImZkYN6lFokRtul
/5bhrMm044jhu2U8jBdVz7343o2gvoTo82KDCxuNBItmahLjnlxYhuQ3XHqkkP1LBwwpc3nGEPs6
87HFDk+RxOTTQvqegHyH2Ynhrn60QrFT+wQxARiT/1jCYdfXfEFh9lDb592oUwOhdOSgxJ8NVNVQ
jG8GpbuG9ZajCyKC0WyM8tbVEadNNzq4GyGOBU/BJP2Fz0R9BVupgXNkrrR1CXTb6E+u0FMHmC9R
YKm0bZtL+sNlqiRD8plmZ7807XimE8kQ1doy5I3Hk0P2c9uE0wjnmI6BVbteS2g3j0gGCUktRsGK
TbgD+YS4bInUfg+xrUgcT1A5L+aV9OnxkBOpHp+/sl0lhUkl8770FnFegmd0eOkBIV+Qx4F8SyDC
mYHrzJVOnozim7/CV1NOLuubtx202Buqsl+9nh0Hyj5FDonTmArkdozlVZK541v0FQQMJ/P+iwd1
KQCPLg8GtWiHhtajrJhs8CL0rpcSYLPuasY5HA52zJmOQ3BULCPqyCKLkQsxMw1o6XNRytSHd5o+
h0W2MvnDblotYp5i6rLlpkFYjgNk3us+NmK0C9p+2gzRUQRcgTHWJTJRvzkNkq+WTkyDnM5vJt9e
jmKGnFnn51tGWxcCCtP4sD4bX1mJeg9vcuKWoFjnSULflbSjebQln1ret5M3orTS4zTZXmUjPRU5
+SDMXLzwgVDNCRJBBt1s51dw4NnmoWKE7nGFWMTI965WcAme1ONL0qePjun0H8bvIKufB5lp3I6D
R66hFLjNDu8Pa3h/BgJf3k4Loz7EnAFBXCA7YYfYeVi/gl16IekSGBhROh27I+6z2H2GESkmhZz+
JXBn0R5b8OH16bdZUnkhFlTQ+YalzJmd4sLFBBP8FY3av9rNJYCypHWfzax7VoZHPfQ07MIJKJdi
8gHLMYUHybvN9V1F9TNlHqV4/eqGPDITVKM3WSlZlRMQxmQpmD+JDSk1je+KkDtJyAjKYJ3uoVeH
w3cUr7HY2CFO/iwadkAdL8XU+/3GW9AbDI3SEmXhvCXkH9K2N2upwx+fWmAzD5cFLauxdgnHbwv7
fkl2jg70gMQBGh5vgrbadAYoaE9v6rgaPoxQ2Nyw6donFxYfnvf5fIUtAyVSWBhlq3ilbG4itoMv
JfNDm9779u1thQy+7RBEo8YHrOCkuYhQDD2xu89eBpDes2n4sVQGo6sUbbKsxXpSEU+zh5Gv2Q8G
y2YxEzgOUqw2CxevQ8t9kn8aY/374UsMOnyqUlHaw75OTXfw1xKH4azjwV3tv4ZV3nIy/7FnT43a
td117G/EJR8nySLtigPJhOGC5eh+fEyxODvcQ7lSGE2aw/Nv37iR1Tj3yhIi5quXq+bw8eb3g0PP
L9W5cpE9q5SQD5cqvPVEguzUAzcWWuUfPTkGymZupYIviPOf4cJXT0LP7h7mQAw2Zypb1uZi5P01
oa83FwA3Dg5NCqbT493XzQ7Y6TK/QEAlRlOF6JHkMVwRVj6uqaaneeI8XE3eXrrhwGahWb+foVfs
+qDD0RhQnzVfcxcQY3mKN8fI3gbTcL8ad1GSqdXseMUVg/MTd/0ph/9Sb/ESKnTEJu/tXVHpJb5S
HR07HsWzby6xiZEhcmuAzLuIYOSdRYjLQl1COD9JV2e0MvZciNSXDoBLe75R2xeTRvJj7cTFvzPh
8MZE0vuopqmMWb39vuvs5/IgBGu5GF8tzmyi9y7Z0F2tljYAW3rmSuukJolBqhpS4j2CbxXxttvu
FNHdRRcMS5gqRBqA81SguVcaz/Z8RjUEhXcZ7DKfUABo4oJo4/sagFc1OlYhyi3mL9fP+CisJJfT
F4jD9smsZ4WvVqIF2lURxilYuR+KQciX5s4U+SCAOHsodZ52TBIwKbhOao+EknDobUWjxdce6c3H
EYa8NOGWz1SInYU/sjEj1oWYlJQd8RtZB2J14ovWCW1jyMqG6vE7mZB0Dp6dmQWsDPF5Qx8oAyso
SifPOe/yJjGOBDVjslGWwoVeBsZ04jizGOPBCeg7mGmjWIiuSWYfC20C8gFieckDiljQF+pda4gk
JDwZDDQLDBu6A4g0YcK+7XKRLEY0n+88YbmyTjHFGzaQt+Ej22QbqfbVEdKKdgzIVhRTFpGiuYiz
0ZGnMdYIn82J9xB3yq3f113BzTJwY1O8gFC/aY/6y9FZB9z5ngK0IfqbfyzHTBKL7m5ZP5xYcdwc
Qf/StYslCjkWzJMe9sLrwPg7mAZ6+PzJtVs9mGxbNpXn06Nd7TpaxzmwUsKBv4S8RqdMpX5gjtVT
/uhfGbeybFV8FjffTac59s0Ftj2b6wz43a9efxdP5ZKDXP27P7xtANRZJEs2bBwlnWaedytDfFsz
reX3Hi6lTXwHMeHJQD5sby9VDyvL1SDIF/rE+pyPRLoeFH7F/g9jfcSw8pXwKVA4tGS/WTvYRT7K
eSQO3xaNrczfynehV7hS2kUX8gu5QBNFTbspiyzpIsusi0isTEH7ZWOjnrCzeMFSHCy3uox8kvgF
VgnLFRv5Zd8UkSrQZffWHWiKwENE8ZIHEl1WiQ/abSKtIt21h6TZy1axMTammMjSHd/k1DLtjSgS
UbDzC5RdguehjygO9QFCwSAR3nf+EI6ggE5ax4azJKoB/hJhcGogIFr11pc3oJYyHWGi1Ykb6lQD
ndl1+RPchRy5NHAemUVBt/Mhu+/BSD35MMEi7BKbN/BZWE6Ej0jrYdtUjpqZiMAIEXSurNyJj6ft
GvJbrXNL7u3Fgr4Hn5te+i/GhGF5NPf4HOeRCNAxbHaSJ11cFHNSqmJUYEiP3qWeqEHseiiZHw9r
PdIs4fh6l7QNUlOXqOjxU0DVAkdUN6K3Ax4U4IyXw/pKGsg6C5gJCW3E9mrigyW+s9Xr5fWYSZXs
xVePRYV7ueKA3oFZhUGxmGFLO51ieS/GkGPXitaC8I7xlq5t8tOShfGyOswVIk1iCo3P7pvCY/tH
S/hKuwjGjGplKBPCB8IZ9XWoxTo1/UBIMS29fOXvul7TcFiIifD0KQ6Y+yp+w1npZAWc6EWT8gjS
HkiWWQu490/EKcDpeS00UsAm83rD3h7sh7NylqsvBnipmUztfFbkFBtzPvbK8/S6JdCDeBBd/Ncw
xGEPC0LsLBaI3Tj6saoTvG5amT0dZxyibtFKzc8LBb+scNGpdnmEsqkPLBsZTXGQfJcAq50m6BIs
sjgSKLB/uEVWzczV7/wIRFa/GnU7QmD6M3bDkCnWVs1ASnmEFiEHpNA6P6OFO2XCcDTHB15oEhWk
sxqtQ5YaDGC/FF8BgfOr73n+ZgLBCDLa63/M4BQfN/Qj1kaQzGUHNND3Y9hDVKlcqsqiviElluQr
XEnwUwQ17jjdZEQNEE1ZzuiYE9lbTx3kMNI4QGT4uboqN3MfyZP0am5NPzkK5Li+WLFPIVXw9eu2
++sufK7J4VvjYEZ8RCY341p9sfkeC2/tBaJGMtASB6uaVpusyUkRKBCuMi9GQjnHf5w6fpka/h/3
w4oeCebbW0bOY/PJBhc2mJiYD5CYPhLhyHmkV2kfvNDCE0n0Xh0lkCnajAz06ldXhoqmOyOnPq1s
t7uPcLLRq1TzNQBfJp0gxR2i24Rc/Yj2AicstloUg9iD5/Z84oEf8Yq9Ierj4nwfq+/nCbw5g1lB
CE5z3IjckG1gFkMN4WwTVkyms3XOpElGtRS/iyxHPTWQqo2JlDrI2mrDplPCyksH1Y0W1rj3487G
E1VyMBL1wGZ3DMxYq6C92PSc2Cy8wTOu2T6GTL8K67GsN7W+cHb9fRPyZEzST4jWP7FEENSjSvlP
cwXgKWYIMrmgSBupJt5R7QY7mQu/R3GkTW9FXCMXb/ax+YZVhF9a2ChhrxQYKh3YfG0lytsxNP2T
GWEJE/D2UQMBGQYm6oyjz8NQEn3nxmFcODIiOl8NRkjz2B62UOlsMpFHf4xiXeFuT+g0ivsnoPqM
j89vi7gHTMMpfo5hojsJ9FJaK9s5Gg1PU+Q9SMzqo/4V94ZWTx4MWqP98ljKt+6pGBhUq8lSvq4q
81m4ctASwLrqquJMHcBGwY0NFh1Zgv+R4Urd07vUQmSoLHifh5+VyjEftcpzzaBnHdQoYCxCkpvX
YMse70PKMQd9MvVyWwgR/6RUCdj1itbrHoqgqCU4B8umuInmXcxddYhG2Bm/V37ZXn2UOtXBJple
ZjTCNZ3irTy7ME6sWBYFLeWJtj7ZhFpDaE7+RrW2U519F4dWv37fXtjBi7j0STjW72SMYdZIDR55
O+NpfKL0yRuy9577tSXP7djc3gg6SYTd07M6TEup1l9/m1HbAg+Uq7TMIizoGeh5XH1cHYpixGOp
lqewmMN05C/qjdgv2JcZcYXcswoSY7A6lPN1mXEpwWiv84yJyuxfna5M83AV5nbN70Bv8cp0+vKl
plxcIo0bv/vJtblrsvdz/eUQa0fP2twAqpMlaem2mGokipbH/KsKtaPj5hpv6hfr8kvsHx1vls6e
mj5xayvo2cxZjV6ZRkiZSA2FnLBzYU4f4KweM9rSgFbbpy9nXsNmZoVLrTQYUxbtFXJZUI8YNJ7D
5T5G1PbphkeiFsIJU6XoaszZdyyej8eidJakkLGZHra0pP73ZqH4d6p09mX38hA3F9XQKmejuArz
MVAX5preRfYHNVtIOyhYmxyqOXkQo/cWcl4WsxtCiT3I6Bw2sYx/PJoexVNbcFclc3imMm0RLCCZ
d+u9Q2+nG2IeipYqUZ79daOJPRlClmQcm5kw3uhYBwch4nnoyCXacOHAOviro1k4P/jDH7Xps2OT
VP+wMwENieM8kWkOZ/fzRDfGsVzFRLAJJtlYh6ByV7cnvap89+lzReLJO4lw2SPn4+O6vcIk2tyD
dYLa2tilHYWZ3EkScMqxUaWv1yw2IsvmMrjbuWIQbSnZZEb1Li/eSqjARo/FFwG+ETIGvWsVqFA5
3I3wI/8DZjdiSUZOLTOm7Nqlec9TI2LQSK+aBNjUP36Haw1t5jjpFbekExStjQwp0gUqwm5JuUKU
4yNTGiYR6PoONXavAnJhBiFpy4o+Y1Ii3fJhSK41gy5IgIylD0CHMA04Lk2F3d8gKvEYma8cSK8y
udRnMuSTfQNl0TlHgNQ1rrASrRcPFsbInyLBBIMQZyoy1y9asb4cAsCpsvHDGVMcyOwwlEM8dNuY
kNRdtv2MoXCV+7OYzHrCO3JsV2nAf9RKrNbsPCdBiDKmZJMH03KIdrrTss1eGcYlvZHGDZVw+d2P
l25agCt2zQDR/Q2B72qaXS/uT/lqrnkMGSdw8denHHpA4I9B9uOaLoFknmdFDI5InzMClsLA1uXf
S0XA1jzCqRX6oQkbAVyAyvHrUkmj9km4F4MLZEJKyGIHUTGdLAnxC9ASetS/O/OXUdKQqCB0hYCE
Up0UEaMLhJFe/O9ep0YJODz6DzmLHGDoWi9h76eZ1tpWPLWcQUdu1255pylGZGnabJr0Wpy5vO83
F3rm5fGf2KcvH+aNxfU0fYV24+EnfA3ffJWHSKKsvev+jye1LrIsGIRvfMwT3QKscsVTi+dwpRzy
pw7FeIRHai+ItVAEra/GpDB6yA86mbdMjaJPUoUTd8KBGNloC6Co4JYRwlFtnMZDxxyZwflxeJBq
ps7y9W4yDMBkavTdIgJNNgcEOCpVVyV7aVFKN4xxuhLdZljMFFt81tipEDdJkS44EUGm+lUAgezH
SYCiBvBilDWzjnms2Z03bRhxy9NISwXIps9MJcQ6dXMgRhFuwg5GWGcS9YboPsQJIndN25yWuKiO
lmmYBH27SWJoN6fnrFVan8OV0TUFPHVDpvMaGFXNkPxZfH4dyNYIEiRv6HYHA0nwgJr/rxthbNSj
otTfJL0+OmSrysLG9kGOYnEbGx/SEK2toltxyc0aopHji3XofgVdlNvW5a/9e58U0yiRF0gEKNcN
+YrEWM7+A6l+a0n52FqL44hgmgHZ9w7pX26waYIA62CDOXGg9HdFMVwNwilOCdFmCy0cuoI5m8Yh
lY38rnxaV6olRfsXqvzvZJy1Xbb4nEQo1mnUywXnbfg8wEniYWLSZDsTTRyTPuN7Mrt0G1VyDCZk
jVRqIrv+a/te+/nFwqr0otWvpyS2lYytD/IzVtWu4L0qaff/MhReHJi2XLvYTv0dMZsFyvPYmhFI
OHIqPa7d/iUJXJgU0dpLkGouHH3WvrDNQFNx00HO3n/ZnguImAY+bFvF4j4W9Qbj1L0Ao1jlSgmc
mC8z6qQ0XWxkCKHMRTGE3NQ80kxpyEIuASeAZz3KV0Hy/0zu3bW/cwvIbJ03b+Mocy77sWPatDaS
dZBl0t+GhRUgN5Edu1P+vFrRuhSP1qxSlQZxH1cuhL3uOQeX8Xc9onCKUEDrNPUJabGbKKnA48Q+
X6gWuEfVHZXks5xErWbBHgvQuEHATX3IeArFyOs8g21y+FF/7GrgGqro8sKcv96kUZzeuUQg7A+l
Qqr2iJcGy9paHJMl23Mn1/630nfe948gsrWO3GtwmFHdLDYZfpphoxP9KS3XorhQ50HYbjiT5LaF
SBkdhsKssM1kFnv5BV2c9LPpePnmywgfMV7wPdQQlWkbA0x6VoQvcPmdTdtWj55h8CJlST4Ac15c
SPT4wtsYgJZIDnMi7xDkmM2vq79ciGWT5zd6FLA664aj4s/cBHRweQRoO+IAVxJfwfEjSSVqOkTZ
K6AizhMaLDAann+IlImXkvj5xNnBlI8+1RPQM+ICjOosb7W98kiFGMa9jNWV5eqx71R4sXf362I2
fX4pYai2vPAE0FHXCM/rurWiqY9IzcKx702mqsBfS/y/j1UtZo6TrOry2O7ikdwEMOV/w6phJKQF
WUz34JiuNLkOze9IpSiaFFIGZShYm7b7fAhVPb7t/77cXYyJxEhThxPZDA+bpU62XQUYLQ8SqISG
1iQ4DARCpdBTzqKAIMrLZe+kci7sZDmGZLizw1ovVoB4bnxKp6Zkos7+fNgb9/0pMecXgYto4pho
1n+DCtBs88P58KxcAMBrGrqJeKz+xso8JlDhCkQYellfi8jG6vrs86f9mF4RgjrNRo2OO8YTmCbs
AGccURJrGZJSt5r8yNhsJeH2hxfwJwrL+IKoGGXhDTMXwuFdf3ESBJ0xDhhTPZ4jtSKOEAN+xBJa
qlKYQnG3zS6F4ptmYORdmxqIa1IKjAi3Fj7b3dJswHfaEbWGNxO5ZNj8O/CisajlrlQsww7TL3e1
XoBX77Zk1E4xpd6pM+4Xsdbf0cMqOOAvghQWgMR+M+Jt8+It2k4RKXSCEuVJzd8TeV6FFe2LTetm
qzFH9awCMEtYRe1qGyO/e996hCUkkK+f2MamzMLm4lavSf+kC7yMwSmjJKVSeoMVCoNXZESrE2uM
00Rr6hVdbb142CFGu1G1AykD+YnWqFMLCcdeiirr3UPMoKjpIek9FkNvQ/d9INrM9ATGKSMkWhZc
txJWaktaW5XpF//OBtpVZ3odguaWZSlktoWmAH7Ap5bkavql/osJIIwH0qrlJwyJfRjBRJR/R/3S
PHQxNYE6xRHJwLUq2fM+FTPpvxO4TwT2uu4P6JubsTBGqZeyOvv/TQ7dXz7Bo48ppmn5VRsY59Y9
s+hTxvy2MnIm8fqbLzKQnt35D4hF8jr9xg7JEIzPlRNFm9qL0in0C/akNvj/yWLYu93PF0zvHhG5
JLYcIRwRWmRx8bgyYYe8n1FKcCumClY4Cz1Lk9n9bUDqNU3dKnVuyKTAaxfUU4I58UlMQ0ZAn7Oh
iTL794Gby5Hch72Q3LN2VzVBYrZbuexcQPxbIXSCkr3qKzFHNRBbxoRFkX4peURByezVnrVScMvM
cUgjt77AFBtZ5ltoTeX78Ib7ucyrGyNj4+aIvmlT0Uk73jq80pVSmnaVcgug3tifGc4B1AkuAqkx
Vjec8gD8H9WfVE34BF085sRgz6i6K+szG4FzGR1x1R+XhH8IPeE/79dw/rYkq4kf2/6GdXyTthwM
HQ7vUO2pdDxca7tDYBbjmyI5UPmzhEydxcT5i+FRYRcGe3GxSlbVPl5lW6o242JkKNsj+l4EYoQ2
5BENYQkE8Tlb9JcRlJDRYJF6SrzcGaln7iQQ+DYvhZdWhn3oO9U2jdoYVKXrBMrYSPth3GkADAMD
Pt/Jdm5DXeMjY2DI+ewY4I6NeVno+Llg4VZk8vUpM7B6MHwjmxe9XFUbzccXYusdQooFaPrPLFNk
rKHA49Lhm+4sobgrYmq3WO7aQeOH5GG5G2xLt/mE6tzIZaROGockn5++BZiD/BX5qqeNEFw6lvM0
P6UlkkKrkjbKVhxeiabhAf3cW1FbE+MfHX3A9VoAOEnvRHPJ/ZGRoMx2MrJghUoBFkuB3QF5sNKV
4uaNfr/RBx7isV3KO7Y9CF3yBHUHEyweLeNV4+Xba4WCR41MFJi6sSBADbJmSJBkX3jsv7yJ9r+i
0pwIbWwF1leawJNLQr6dnMSytBf7yxtCacNMEkGlM43ktMch4L1n8zFemEKFXIo6YvK+PaErViTv
+KSXh1SLgfGlh8BUbviRo8fb7bxabhDwHhs0HVJ2iAFy2GgTAcdBLiE6nQ0KqiUTgzKywWnrUpHe
QxGJoQIjPmlPKjcbcPfO8HueJ6VjSPRSpsWGy58evJC6Kw67mGm/eNGMSVLWrzClvNseKOqy8xXQ
ptns1kktA9Zfbm4AOdyFi3YcATp4exVCbTYgWCRpyLqhIUJQWS1HAebcMjc+O9huSOwGL3ptMgzE
TZqVuo6w3iFwyIiXN5nxQ8G8VEEAIMB0xE1C8eqM52rfrmaIT9OsuCabQLmKGCk0no/40mo/BX0j
QpzVKJxVr4hAXmOe1MHWze1YthC95xjjUFf7aMkxfmc0CxrwdlpFWXLsTFKcKgmCZ+ys02i+HwNk
jdvKMilxYzfweIFau3kv86MG0VKoB8xb1Wm8F9OmbzPQlMlwcoLzPXvFU/pO0p7zWR3Kk7vpmoh3
+5F1znP+xcfMosS5FzJEzDPUhMH1mY+VgNBVtgA7QdqckDvLN6rcNlP6mUqpNLASMCVkO6oleiFa
njpuRtUjD0UsaBicfOUqd5QZ5NdrJR/b79x6ZRh35Rxv8mYDQDmcRcqDf1G6g7862Pyy634pZPz/
MhQjTvao1jSXKaJ8inO+zgoHmiH+rAD6mb/0W+W5lknvT8NeYUXGefEwxCJlAr8k0xse2vHoxSA1
rboagiJY5gVgA1cJH8CeM83he9oF5bEW+iQEmeQvoFGfAj67FMb7gc7EdZmyfAxaOFxzekrr97yr
mz4u91xq+1os9rcU5a4Oq3q57jxy9moaE3Qah7qdNBjFxJV9GRcSPjDwReRUG7KUIrvaTxuV8Y0I
n356oMnQSJaAfDWdQ/u5TqEczSJlo7gRMo8P0fG3eLUR/HJ0XFxkUtj5OxXUR96IB11G+E2CB4sT
nMJMVmaaWPLhLZ0DjhElWOT851GnqpNo4HTK6vnofrWluL/I5J0gdX+q8dkHOJEH8mg6ybL/TbJ4
JAjje2KlLh4VggezvP5am21C14/OSGzssK8w7KrOYXd8csiq2OJim3pEMWZGuHy16xnvYTpMTsuQ
MlENi+bzR3YexZqsrgiZwZaS20Cz8C5hvE3N56XW4RhSDiE4ER926o44z6KdB7hStsHEmX0L81Y6
vPsoa6Wl8Vbt1eSubJRra8lq4/oI39JHh3TqGeFdZGtH47ARJsvrQr8L0GVI8TytaspgZodEyoZz
TORaMsaSphV1cx+CurTiNNmDVJ+ketn7rAXjYdJD25vZDHLR+3XxYOCvpI3Y7rCuKfIWaLBEy7aO
bUX6Ku64TT42REZvbNaH4kkVGIioCotD9nSm2jn9sEclih2SAAvv3oboXY/29GuOWfCuI0DacaqF
VorsMUYGRav4TRiiGlFynLa53i6IYp4vrNhldvmocOKSf//GpDTjuEuULENd4aA8H9hNljMbQPV5
JSuKOk6XNXX1CDFnznlO8frn29/pXWVW4XFyQZXLhEO91/KsNIIDcW+4w7LTwJmUtbYrniC13uer
QIyPAZ63wmquecpjk+vVq1fOmrMVN5ks8jloBt25lGFULTgpdwCQxtjWPNnyTSVHLMpVulJ+HRat
zEPEsDM+j9lET7nlGtKvTiF4gCXK5GwORTSw/yBFkjdSbhbe9nLpxqx+ncQvmw9T0E8lwgBelIKr
5Q7NzHDCQVsrYk9VcOhElfQzG7NIys0T8lc1HQxBiSRvWxgWmdbcruq2q6UZT6Lwd5zYchDUKnFw
u4ViukPSta9bdO4SP4s6eBDeTj5YATJJ+JbHhcZrsTVz0NkxlAoZ87IfL/vYfZh+8CTl18ADmEAF
8ykBLycxYDT7wavHjk0mdlatUSOVtnUl+/bQNytAstuOLh8EbIbwgqu6k4hFx8D7EXQoVyR6dXTl
eqPGYgyLDHh/Y30jspDuL3tV92FejY2mbqMDNnhZG4VRHet8BU9IA4h4fY01lee8wB6Td6mS67B2
QQpGBVSJTSWPcMOJ9WlRgEi6+GQO/5NlP3CbGtkYlRUKDBXnvFidGUG30XNFXiwivkdQCX8eYj7U
bKYhm1r09LzZbdaU3YfmIx0oHWlebKQrfK6sJm0zdWjjLCN/7Zi+A7/wWpXRnZskKUZ0kybeBiRP
iC1tsXEOmqfzxwsPKWldVeOVzJxlKM/KNkuemoOY9CDXoD4QNMq+LrgfRmhOwD+N/2IVGd6qtQ/4
zEJJg1bq6/DH0goXymLXGSLnhW15unFZRCSBj0GUls77JnQ/jLMhKNkasEwbsG2KCoHazJzezxoa
J0rvN8ixTQst7akscMDf8kgCjnyJPuLDMbqYDVQturb6ykrtQRDpAqhyYeImuFbZ3rawy/h9HX4Z
1IFxedeJjvYkuNTUF+4HU8ON6FljEVmZitJ82VnJRVspcusb7JgPE+LZpgWfnFhOJnf1NTU2isCh
3pRFzEdOPT/sHjskXIu1TXZ3sebS4V9o69edJSx8CqWS4L3mz/lHmt9+rz51PN7V4Fa3QhqvLpaV
srVhZcagu8XlFzdRR+iaIRicnJ9sSY1a+Qb7SWhHxmrUmv+w6x7NnXJ0JUZu5V2rm1CMOQIuCNWt
WsaVbPT9sKYh71Em9hKSmeUXL40tJlhZ030dT9AW7sgJ0VM55rFLfws5x/kTh9XeZDrLwgLZW5hv
55tqUo1rWAy4z9AK5wmx5yvZmkgchvh99cPlyVpiHSJZ71v6cA967dxmI+3ogk8m4UNjYe6P8sA9
db0QuihcxevsMgdvubco+OsJ3O48VuMihx+Nh+zzPLKGPDjh/otCcn5eDGa+YTm/ZyPu25Fd6ul0
WZnJ6wypDAbTxS//3k95u+5qmxt+F06SvdY8/IokGbECReHZvsTaa96rgA02DzXNPf71lBBXQ5QE
I8AHE3Uw0DBAg3EuWM0VvJ0Q4Z8zjl9xKxH64PsT0CwXHlT0BWoDEEHc6Qvv2NsmYK2YFUM/HASl
ErWQSyOCHMaPjqoslwgQccxB2QMRQcmMSuoQ2SPQJp90RF+thk6rH9zbXjQEMPERFTjGoA4U1bUH
w6rOU1daAke7SETAXSCsMcvA3pbQXFU4MMR4aKMWE+//m/N+eC+sN93ezCPj9W4/d36qnP4rJLfs
KyN+zk9R0mpEkFpD+X7hS9yAItPUCZ5UBhHjs/N8vCW+6H3FZLE1lHjryhs/6ILB2XrRLGIUOi5+
zrs5kWo87euHfnJJttNuY9ktTg1DsGPTcSKk76YvH6+0/FhEN4ByXFc5JlnbKg7pTwjfjCj7IEGN
kf1xRWULzAvcpqJ35xaODrVFdcBWdyARe7Hk2qqdqRgD7/IOB48IkoANF773Rm0q6FeJdkNxLZHR
WoBgTPCN9lP1wjAEo1ufpmevuEXdmloZ8zeFqUKQtanyP9IQAFeSR23PlP10Dd7IRBMMvGU891J4
bLuQaL728trViz/wX/G1sqTnXF8qPpg/NB9QMtGjVzPwC2Ma2RYsiDkCpwu4HNbQuGKEktJk1akk
pJUoPSuBMMQJWwF/l+mlpVQL1VZrdzi3IGe3U3qr+EU054UdP80QPsEHv1g3w8jtAWJIwimo6wQr
9BhxUaxntzz04J79+YcgHHLR7p7qh1iwbtU4OkBVoAxsxK2LqeXQvmMMfhNnJlDrmnjhzCjZUbN6
34DcmEVPkHOw25zCTt9ZCgEf4S2V5YpdgKIN2NCOJPFzoHY9YwPcK7JNNErfrzU6/eegGEV8lCWh
Cbzyhu7Xb0RjARgc2fqaAAaqD1OW9/GfIArfkO/HykIhZ49GEyeMcP7GQFJSMruaoBnoV76eVQ18
yzSCAjcoNUB7Q97b8BfW2AWGU3YFxcmUAMyk7BpGws3zuvnKrnY5ky6fz4eD6V4403Q0yStC3FlG
mMeqiV7UaEHAPn2gguHXaMACJECJVhNtbxgEEeBtqPdsSkVQ2s56Ksx9vCmQ9JVuooZqtTNiGhNs
WNBTDvKwsrgn7GhP+hVg3k9Oht3pRW+3yc/AsVN1EI67K4Dwn5cqUAn6oxl9Ub7V/xlVfm3Xa/e4
EtwRL3I8bZBpzQ4u86XU6JkFwSm9/Uut6cyP/ftsPEibAmbqnmpeaIGmL3MwgZj9AJCavR0fVgzR
NwMuNyi03L0F1LTUfrzGr6YF4476E6n5sz7/B9++WQQ8+X5a6bdmlWxjzzRQYYvCnYrOxjuE0oiL
dw/6m8Lrmsh6u0kTsJ1bFyYmDazZmo+12Gw6AF22zcz2tuF+pWrXQUXUO+JlK7qUUKCLHOSYeTQI
rmLITrzYSMwLLFta0zShLK0BqunfODRZEZtZ12pt+EgxwI4KxhJwAz5v9w8wB9fCcPmT2Mqo9w7+
BxfNrE6WmvIdZICtXnsqys7akI8tdLcDPcJ/ua2vliUAhMvio8WTHsicmWH09KUm99Db/mkj6SrO
1Q3FqZGjVuVWHf2YWQ+Yu8uoo7RwIOhCBJJJY3gR6NEGiR7YCupTorguVr8ZhERkf2RDNIKN5AlW
ZcwZj8xZaUNlzu6c375utnGBq2YZ/5ZGNDr3/OvOIoxSPx8ySyJwu/YW59zdUrrzOIV5ZZbZ28RM
BAh/M5u2pdy8DlVaSI7/vTKWoQEuVskkEalDoqfvAogz5ahPoKALt1I0/kHUJfFgVHMh+IkZSucq
1KsSWxujQfvx9m6PR/4kDRzc/Y0k+mE84Zi7L0lzxa5NDPjdiA7Oq3ZgFyvx4niD3ISYxaL+DuNf
ZGIVl6y6vyH5kyzE61LINCnFVphr039idKtxONZgtLAHhA05UlPepiS/f4oMsHnOlGwCKQMd0T5i
9zKcHwZq6CE+mUNkAIhz6BesqsZCA+QHAElRs55Di2xk/rlIyzcvnBHAVGExcJL5hyup7KL/pk+z
4Ef5wFuZMeuY1FpsJZrn1X1A45/ERrmE+tput600pHicdbnRm/GQ8kBSYADmyPfFNyKNu7YJQnGe
YYS/VrY47Y8wo+jWaClpWYaEs/Vj16GY1zTz8HBqOEQSVnrR7ZtQXKof2MK/gSkXI1jk81Er5VXr
l3mymNk7AmIO6UGjYgCCR5nDweI2MaFRj6YS/w91R0W03nuKcJtOpsKJNGDnCej+2ifrMEY0KOTL
+cAfrGEPCjZSciAFgsIiDycCvzluPeoVrjPrPL07Wg6CC1EyBib0lhh8Bt/FGhzE4oknT5BVur5A
4E3Y5ctTVaJ6ysBvOxwwR8HORd9QAiWJQCblopdKfZIURBBwvqj3sI3QPbCwEf0Uu2NdJ+upa5vy
TD/vqguovCyiZDz+ewuO8iCKF0ruy9EwVi1ixtRtydiWQuusPa8xZ3Li/BTR9pSQrniTm/a5I7yg
usK/0fL4xwVA+8EPeLDqv4FNjoM5xIuHbbvpbU1inQUgLdtWjYCoo95ShznGBlWAIK0F34AU34H3
o/2h2istIO/kQ4Q5KzzYsAmM7GoYAhINOApjPXePlZvqSMuRgJj8pvWe7A8uGxBikYvn1hTp0vub
8Oug8aGVzPspslyvVRztJrr3S+qmMJZftjraPG2hyVPcTiAjBwBy3TfikLOcR0tE6mU7F70nkyop
dk51RU56giV2GFBhk8dScZnBT0bWvJGHB4t7j3yZLFm0Y9Wv2zXayAkXSaJ6c+8EpRHLIF2W7pSx
QNTNCqXPm77QSI6p2YHGQYtpU38lkjbbP04+wuH6/OpqSPzSRY9oPAfLXatlkH7zdVVwQUd7bwkg
3RzCNhuim7Apr+Mm84JppYnZiIhMx3sTZxVQHiicePPKBqWgKS2ovLzdCu2VtrRQf3pBRQ/CmOnh
LVdc70eIsxfhjjBe+QtQevdTj74xfNjUCLVMiZFZbc8aenDh0lQMw3IaP6O1une8wZD6fouC7yQn
OxfQDuD5S3CpYcEcBzdMQUonkViLphHGNo0Bc+bM8uw1nSfQX0K88R1Cd2yWwx16/NpBECAtsOsR
BuF8GBLfQEPmS9aYmKWkj6zT+9e0++PNfuJ7+DxSm4L9W0xWEuVhdugSzpNn0zsqTmeKqxQQ/upq
TUbwTyaoH7xF5Qm6hNLjwDCo7Q5SyT9reb0sZYl4RFDJS0U1dxp4hHJ3YznwcXgi/S8Ho4Qe1EOh
wOu2kEmmMYdszjH+sQ4rrLbnVM8PYmKUjdZBvVF99OZdoskF/a0qo4xA6TbsobBSsQAe/PTsUnET
N6Upbk7Lm+3BV5ecDK/S+gx/qoAsMpKEtUy9cts9346gGTAYrghuYu701onlAizeGOUCqZrR9o9a
HeaBl1aa1/vCdndPWpPiXH32xq/klKNvQAZrKkT2Vd3KnHq5KOckmu5rHp4lb+rRldhrLU+MZGQQ
1l3zzYKkJ0jrXNyhYLPh86Qw1fGC6JgFkMzMgS8X5kuGGtRSUgJROk+Au0nFLgIHAYnv4YSJKNIA
FN9AU/1QJtGaP5yfWdOX7GkE6PjzomAEyd/hzx9i0QDXiSkxjc94TkVALmsTVMugF+X5A3SYgpIn
THts58eSGHzBidJEAzQlz/tJjbEYiBuzX+DFiXv2VN7qTPl9Byhi2MGqGTlZEnS7g763m88t/csn
CbfYacHQyCGfVdv9OgRUdGRI3We0xoZ5l3V6QGtDy0FVSrseLkWnsmVc92h136ka4+o481yOWjl/
pwdifJV+uYTRlZef7S5PFj7MxHF0VjxJG121O8DzXJGy1VhCnLSqmC4+Fi2vNcJgxsbdW6wQOE1z
wAc6kd/Txo9cTETtGxG9X4IpkPX5biTvbug4vKJkfIIPSDrSKz0hmF6eTTQacrRs7hSfrkXutsVn
OyHU2UgXCBRlOqXJLRpQwrKLluNL7HXcIMNvbwwkfErGEe/XVdCT4ANJsKf99AuqLUXPr6SAF77P
cxi1YEzoaVJ7qUpXae30uvnTO//Wz49WRVo2pJboWVoP7UwE8M2bV86J+l39J9cC6CkDm2eTQEsR
MSNpX4jQz4ECPgHdOQntKrt9Nk938/PgON2lKcYDf9P5CP5A+Y5PcMx/Y+umQ46jnoxG1fRsvTyc
GiSo6GqreJEsO3W9jk0Lm6aNNNmoTpfNUQqDs83uDI+vTSPi5yiEGjYeRc9flbDqQ1p+YvxU9Vqh
uGq1FF6rKEdDRQ4AcNBdNdXbc6917HfNywT7N3KP/3M+mofV1nt5eENr+jGv6MoDLNUGEl4qhbLz
GrjlqHg9TMuge6Q33OfaN1vZ999q5aN37Y2ulXjMdZc8s8ZLMr1elP7zNzNs4I21qf8jGdcqfUXz
GWBIujs2LrGbJeZpScGpQrTeWY7MtRMyhPw5mQZWOFhm52+NfRPsnaQTb1ZInagMhFoYgu8ip3sX
iXZPZdynfIycPAZO3+jz2WfMFu3wlDBHtPEkZ4zhJU1VqwAu+xLME36wBujQZa+wCBH10v4xyL8A
tFlARKNAEJWJCZg4tA6oWIZss+o/VTz8A0kXaUR0bO6cbt/aZbM4p4zF+ZIq20TIch+F3y2oZW0B
/NVS5bWMFINKXhQR0VYlPp7g+e0L4HwlH5f2KzVlCgPoJZXafMWIaaVDrZZcf8uiG80r4Z+7VMaW
ArE0PaQqxfH1p9sRgnd0BQO3gDBGBoB1g587kY4NauZP6kIUIijgLTiauzM08XywnKdiGX2HNh8b
WLhd7W6nwa2qQikHemOykLgCG4vA4i3DRZwIEQg89yJFErVOQPWeqMpGjxce1dzeZWMmXPLVh1BF
z/WgY1IGXlQeE5PpbRn7OyTccqUzBCzvDj8dX256draNcJmPTJ7ABAnkScr8h0XWwGDFaSZ2rbnY
8i2RIta+F/W9E2jsBWPL9G6Vz1JNS7evdCZ8I8icA0PaWprRVehDzJJhCdHjXxhd7z38Thc4j20h
0471sxEhm5pEXjiOt4thA+8k0M0/kQizkyIZlIVXeHc54DTzI0phfemcyr2zNasOOQImmHnBNmtu
utn+tAj3TLqpbVHeZqGJ3VpOWyEakBT4pxBnHdTpEbuz0ULD0E+ua1iwiNCRC63ujaeYMVEJfV38
0BI5kFwQiNTHhHBn+hTx+SSyonnPiS2xF3UMUYeuOh+6NQD8gMnZBTa986Tvkvk6q0zkOrrJZh4h
Vbyf5liFMJm2uDGCjXTzS/NONwhIereGLnfMdKh7c0kgh/P02o/H3UtW5mdnBjDjuOf8qXch6Fpe
L4XJxd2BENTPvmlUItuig9jtSEwitM7JJUhP1g//OYJCQewaDkKc/Mp0c6d2xdm0djCtCEKPHlzA
rnoiaj3k7Mado+zQyZnFt5nwZKa95wo9jXU9zJlu2yIhYRW5vU0KZdevpWyZTNiBYfINMy/ooljp
4EUT75TNKLzr2/uTzhD+InzWpQ64eWkNokjBRNIJ2eN5Ut4PfA0jLcerpGF5g1WL8uZfMdKhHoK+
Wm5Uf7Zz8q0WgSUDMGDe9RPmdehck5WBk2q6ClpqC1CL1wD+h4wsGT964a/ESub2nPYLWA+i62yo
qZypVGyt8sDsDoi7ZyX9hSsmuuwOuC+Bz0ghMgRjLHn3xtw4JF7ppkL4t0qNcV9LIAlVrbMiEsVg
7Dw9zpQMH5WBJyNBgudSsvpKkIAOcTbigstVuewFQI/t+0+AE74uYPXI6Us0u73EVolhrbKkcUjk
0WDt3j3YzhOtM3+1WW6UrdMRk0PFIkJhBnSBkR5KfXHeTaYFca0Edn3zH41vjdPiYe5nzoMhbGfq
7oOj6eLr39WqYoDpdwG8bqKdRJ2qDTE0MmTag8K1X6TgSCXyuV4oJB9p1RR6u4MMNVWqVZvbRK7W
rqmQn+SyL89h+os1ray+RZHCKLgO4VAwYMQIZhFPIGx15+DMmwu5vLpBeX+htmLb/Kw3ZfgeWGcQ
vE0cw80SnTQy66oozoVUNX8t3MLFV9IIHLCuaE2UCOfA0hsRAmuEY4kHdEs0UfqNm3MDIN8EesFy
NoZatxbx7dvhB0wMr8F56McYJsok73iMpGGJmTEhtIEPIBQZdoCYrHGHyoIOk3+2NVi/6Jzimhe4
vK+3KZb6HkxYR7KnPP+iBfVI5uZ/Tkk+gxM8pWKc7yk9gkFyGJiux0PjJJvXMCfDcj/faCC1J2mz
4iNF6SmwiFUhxSrDwK+JVF+MJCbhpAiG46uHNrkyQ/TL0M6c76QEzQhtitrw6e8/l8HlozDldOP9
h2xBjgz5fP0qmTbLfegDPHHaiUbx08rxuOmpTi+q9IHlDCkQTS5qblYv/Y+4jgecTxAcPr+cBGUw
nk7peJJmeGIV7Y9Mau+SCPyu4IZQSlM7ST70T6LmUBAhLGVBgRFKcTI1RqfDmSxfahMBO7+Abfau
CChcvGOU4OlIQ976tQa6yT7RSZOfAcRbBHcqUF8I5RE1vr5f3BzX+V4oPrfS3Lzcxup2XHRB8oMj
zcm8drmfDOCKrIt9//03GCP5bmSrUhUWykvf6dmzB6k/evYGekx1QPTKFbXt13aE82Dlo4x6cIxL
R3+rUpcE08lk+Ons20cagenmkjDmNdxE/Z7xnir+0f12ujNIs7FSXqy/Mc1jabHriBwdVYCbzSCw
2DDvn9MXSxe1beuVXgg9jCoC/0WBgBretPuM6DORcE6+n4O4WU9uHH5trpZpGCZWh4qTeZZviz3I
hD+IHM6i4FXilC6hAbT+xog/wQ7YzygZzMNFmHhAVgkSWuLKxhnrwVgCa0+86PJltA3UKGQRAD1q
jWeEByaBaq9FyiH8JczJuSlRTXTkSiz+VUVxprlhCe8JKk3uQSxYVtGyui+1ZJtAcTxBEtU2t45a
wqZTH1AnPKMC4EuAezdNzO8c1ahVrx9rZXiWp5z/im34DsnIyl/KUz7PYtODxih/Vo/94OVJZ9wd
VX7+YeBr87qNX0sX1TsVboDsfje2yGPt4kTIoSb9JNJx+W8ntkgwhfE9bgVs03oJ7VviAGgLfx09
QT4ZdeUorSwXqpSqBxn53MzhQBR2x1J0gvzJSLzlvTTmWsLtGVm9w7L8GfmvOH+voXpxXr8pOGNj
t4cDyjrp6H4Smr1wF2sk+mqy0TqboRjUPwVfSOXwjpt98QCzVE7AC6kYNErQiHm+WvVdA+Oh/LrO
r1Iz7O0DYxabEYuCXZAuLoBrSVhFksBB5JA6FtfmjAM6J579wTPAptcY9oauz18J81m2bdKsj2C+
UV+UejuIBpG0K6mFaMIoOsj868IcDPq8aAbeQJv5YPaU9fP8ky6iAADR+UTbntGp1WOK56w6663u
jrHv7jHBwzISrL0NDP1om7z4+YY0t8uP7/xw3gSGL/Hf3sKXCCyKh1Q3T6kEmYm4+O9vBhrBkrI1
iViw0x4Vgu19+WAJFFmb1JE4ymTq5NscTbHYoTWsSQO/6lUzkZhDmSnMcZcHckE8wUZO50L5R5Cd
+NNUZHVPN+cz8sHsa1LAt4JrkrxyJ8GCDaOcTfIBSowGuw2uolaEKjEkXh6hQqM7DtnonWQkelVK
2FA4dRM4VcibEH8ghNBD97RjEASiLLdoDwI39LD3x05e04gbZR/E5hdNozBNQwHsZYRmVHF9rq8/
/mjnjvZGzzlRvFnFKF94mhbKghjLMVFXiBeN0n5VGbVO89npSzBJcgs/OgGZU2dYZubw1wyfLiiX
q6DjcdiYNOAckeiScyMCTEir1Zl++8gAo3OXiP4uTPiPV985/SwWQQoQU8kZgPHj4LJcIrXz7H5k
yKBw0t4O9xd7ias48sVTe1lyPDII/a6V5XUovtKkXKu/7UxKomffJ/bUW3N42s6pBVHl8LPSRjJA
GX+/wbXmFhkF7mywQCWb2UlH1tH2lpQqmM/UdhriaEwreRLM3yGr3r0scJF0yh3Nq6YUn1oBtzgB
m3hQRUiB+yYm2+90bZJGcLREAUVKhj3Ey0mds2wUYDn8UyVGhAOfzJcPr0u7JlEN9Z5iaXZpyoxR
a0K3xiAGbCOY5ZB6MF3wxXJ9fsy8dcdi1igKLLuORCGhy4Qa9Z4VWDu/ZUdaN9Si7noPg4DKa0A+
+Dq0n0ngsagjJFwGqTv0JQxDvDgIRniFL0N2mlB+0vXwpiTQH/ZzCpS6HtPkx8wEpsCsNrCVUBRI
FF6JB5tM3LE7cqXNZY6P/Cxyb5YGPcwZbTIBT0Wobpq+90UowukyDkHYagwRDP2XQexBNisaYwBi
yQmy89VE3gERqfgdbw3Qzy/Rz7rQ924EHHXqYaUHkPsuyA6rRDsHycHms5Xh1QhLiGfOiKFU173D
yio3/AqCfxRzBnh3aRzC/qxGUdSgNYY1tQDp4QQVhiZ+0L2S1m77jJC58q1wjP2PnUKp8ZFu6We4
rKd7ejYkfUpbZgHzzdf3Au37/xN1+p7a3lCPJ1i41CiA2zwWrHupk+D+GFiMo9eSsc2KJY3oBLAx
yHngNhOLT8YvbqohvK1N4wNKz1mV5v9B29B0UiQ9K8q2yT4raED9PAdvajgdy5qJVsGzjpmVCRqk
fE/rBNiimS9OFt+hvloavfXnR7yPBFQNujXc15qUfmrR3D0SooXoVx9VDi0GfWUgoo9aemJ1aEef
FP7vDfOgHOcd5FkJ0Kaa5WNr3i9Afb/sc/qIiNqpQRnvtTKuryfuXcQFL2h2fHWgDvoOElcVR580
ACh1sF3cAVZyUcd64oyV5ATpitryIux8KPi6l160/y2Xc9KDH7DKnGUal36mYUYu52rQh7I/VzGu
82ZBkhtWCZqPZ+GwG3kH+2nWvbzY60VnaC0ypy8tRXX3B5DvoScFbRsGy/QRwP/oascvbwDkUz2Q
QAPJ4oB2Pz2RXSu1ML7lEQZlQsPz02XIJzE4Bn0Cg4zxonLodkKYT6+algHz7XOBAdlzdAfk3ZQQ
WN7/kmhksZ7ZmHTadLcUslNFoq1glbIog30mGhPhRSYNJP9Wm+BtcmMBNrFvGtJxvBwXjzKQLVim
EfNKecYfOHhpqxrp9xGbTUi1GMpN0dlBCYKA4oIpoeWl93dvaSb8LiHzbuAeBSR0ryY2rLQKqO5a
wYTpC0OghB5dpjkxKXw3S+ypfdSLM8t1EAYioNvr4hlhVy/+nFUKLEvvy9y+mYOlaS/X/wFrzrjD
NqrdT3yZ6TldWmL/LZqYs0qVUIVPurUbjKl3tuw/LpROoZ7Ml7XJ6oRvwV3SBCndoBd2+AMpfTUP
L0E/6KEx+jAtPCTMjHkY22OUUJaokWrOsKcGQHz4wQ0POsIoAA/cX3RCfzMfUK/APiBftX7P1wkW
wOqv1edvOBirlsMHHZ98xjlWsuz65W7aSjfXnBhRMothzSJErHklQznS0hWC/29fa1akEeyLPOVB
qgpb4nTloDsCmcMZ20VVpIpSJLAx1Q299en1HVlapjplIipxtIWoF9KZAzqM7rZ31WnPEu2xhIKf
f4q6KSTZHShYtDeDJi+6omBlubSr/ghbQPnbijtE2VzOvO3ifiEMhkNlKaD7HN0qB0Qtz4ao1/QX
lVejKzZCozYHxnf4yWk0OwHbUdmHA3zGq6BgBXlVa/v3Wx+NSJg92MNTYEWku1eQRREl/qsjjgng
LfxiKxPszjV0sDWhFWI/2bUdvb+FpNaSRLfNafKCwP+cgv1UVClcjf9plTWldBYh8ypnOiIC0gDc
5OMIckfB8nIgvulHxPmNQWBvPEPCYYMHiw2N806wRp8O62GyGPxgxDMWRrrKO9akzzjwewVuLeI0
DKNBRBkgC9XYc7Dhx9dSQVM19TTPZJYV2dt01v7J1o7V5tRSqPkrtGRt2OBa7H8dXpSHMoC3Pibd
Xg0LAWDgmdK6SpgW1mGveWPs+3h0O904qALV3KjIAMl3cCN5VDNfvY4yB5kwQ1JHcYLIszb/7y6u
5gGjfoURM53iaoAyBiBCA44HyOy5vRnKtw2JhyFcq+jphkAF8VogXRImaI99e/NX8kGy+bMoF3dF
BdE0sdMSjwgEXAdq4KJDmfh4L0HBEgZWU7xj1+4b+rRRFxuaZCx0QTWLcjsMR3kVCThhRv5jBo8S
f6lUQjC/0a68GpvFidC0L+W0lugEGcDuCQAsWJ4exlh9Cpc/GuXT2PdmRGz3iwCjXWtFIQGCdXOo
iEVc7MBtVPfQWE2L/wJacXHmIRc0RhjYJEdgI+G8UrqgI+iF0/RTEvolU9d6dgQmALakCQtyVCyV
4G8k15lsbVRIRUGYGgd5mBjGzt3afM6p64NpWvPjH325us7XOmegDnCD6m5N0osqmKpU25HlkTEu
NPnKO+hd9hMMYRYnSlg898dOBTo+u/SqMUDUmtB0P5JJSJHf1afXru3pFtHUQMnoovmZYtJenly0
Jo/ultYcHnWF+rGRXD0FUPHURRz6AIEst/UUmOqMGQajMxomL7p9eBBHWkrVSKf/lEepZDuCGNrR
Es4pC8GkLrb5V7QVGC/lulw6OdNuWRnnMDItft24GKxM1X1dtsbumvdIgcjiTg4wcJnb5WxeRx7j
qVdXAxxiXIA6StaN6ckenTcVtp6b3Z/KFzq2Hp+Zy0qr+FrQG3A94M1M6olJ+BIChRXksmLsZKPq
iDXqlUDZMNgJNvTsT7DIzltazd2n3CQlcmh5o2Iv5RSWmzZVdTDzBI+jXY3rCVew2WdX+XVfj5AK
AeE2hxRVqdVzOBegmymM4JU5OLRd1BLU1ajHYwXBGln6cHLxt3s8W+loxejLC7pKSlDT9DOqfAAH
F7TugOIsseWMZFC3t9RYEgSEgaCEL1MFH6kt8uXfV2zA3lV+NgDYSzHP0cbX7KnQz/DxgVsQBSnB
f1kRyAwz0gPjr5/Wp0FQNX0YNvdNMdOwnzk+TCyBSx2nVbEOgoHB3WlJipnlaapWfCsRAtQbeyQH
xTqwphfPaqGtamUT8B37V1ZrzGX3IHC7aHTlZFaq1vLiNArz2wrhCguqDbZrtWwuTkSkVFd4EnPc
G/xQHFkpsCK3vQyr9PgFyQ2vtOL6tsaPkbLDRHrKBpPBHddzWL+rRaX+qZz1KMzZN+E3grGEb/lj
rUfX7kcKSe7e7dq/a5NAsehJtA2iWU4vqoLryx/9GkM4KD3qhtHJF6jEumucH5ig3OE4g6yVp9rJ
RBej9RYi9iZt0t37Gg7RH13Pzj0Z+fyNF03DEHVwB56t7YxXqfx6+D0X9PxtLJra1D9QXhiyJWl1
p1XiVbSmXiPpUAWM+GtLEokbtXuPrfVXysKOP1kyxoaRZTD7PErzfiBCRXlNWvgS4LagHOpRCT9y
nbgE/AV7z5qvFazgGGv1BjOy7iBuKCNiBoKzLzBjTKgimc/twycIR0UW8fh6+fx9pn48/m6dU58r
gt9zUzLbH4JQjzlsii/mExKW1wjOKE2rpyvAGuZfQ5b/9v7ls9mZ7ZQeW2R6xY+or2x90M4DywbU
72VLE6R95NqtKGabQoJA6xljKntMjAxinmRYE8Y07GgGqxE1+UGTAzueu6NPYiOAF83rkKz4exk7
DocUpSiRO5GLwTmokYid4geeqos010F8WIzVdczaO0lewzQmRHvkO2U7awUuvZAS9jPEUNRH2ua8
QdqCOoiKDdOUDeyb6wwvVa1a1L92pbdMqhhikfFi+eLSvSc/FS5r/Xlh0Wm0wJ2SMuvtomWbIALP
7IvqnsvnbA00449lxZb8pTPLrKZa9dSc8pRvWn/0vbha6EXCP370KkLXqfAnzEVDnmJfJZ3ZAIwp
zi/Hcyhpoxvr08GHlT1dyNJRaLjRKe7PIwKrxLRllXud6mU121xQIiwyO0qD3swgNC/NXiCtKnp5
EW3SOeiiCkhZ2n9ZyjVKCAVxQMUSkijS4tVX8wFmeTVlxaBpOJ2YnyXOHEBB9x04IlM5rFqSBz4P
D7nzrN6FXQRhpnCsxh/yhoqC/BJEt25WUXUTRhUxbdOZRs8WpMHX6P487d5aPpv1kqbqSxR/HcEM
bNX8RJExHPvsbTNkiwhF7JkCUWBhq3lUDryQ3spKB5Se1L++P8lnEpqn4bJCMIJ6WHQ5fJtbsx7c
eOxb58xA60iQfRCCXz7CI8VCYYe8r2ZyFH/HmnCk7GDJGAmhFGUBmTvCDPIqmkGS71x7W1bN1LVQ
oKTlvOD7Aeslb15/XqY7eqjclwmUyhjqKLf64gEEsRjWQUWMrSiuNb/WKVqUYpEplIBAJIQYIE1m
Bc0nMZ59NXUMG57RVKzvhVmiYeHcjUEVE3+Lnwq3WqxweYqKAh3OhdH41/LtYwnFySFo5qqkMs3G
ZaV199s4L1NiU3noAtuPLFJndMebfJV75QKWDp7e1TkrN5KooxYs9/SHkSjwpK3+xKvBCBpaff9J
9WBzc9bf2GQmVQbmpoZJkP7u00+3MmKa5Sw7LI/41v0QD69gs27juuVr8VAArvotc/iIYA6JIfEE
Nc260cQeSyY2CDunZyIiHdoENxAzeiheEcxd0yr0EUCnzg0FAAsc93DELS1LhWCIAhRBib7uLtYr
GyQgmFaCKFRrVSOGc4TMdJL9NdyUJEHpAam/BsO9eZNVqDzjf3NqFBms7lkELApamuCCLnMbYcvQ
Qg2ftLKaHnMhMl0Tk7OGebU/exVMDOIdmgx3pTf3gEpn88h4swZp21t6TotXi3mc333T2aXyBHHr
ycYmtE5yflx8c48BRjcbDOchy06b+jdzk/g/6xtPwppwEWXb+BTsEpSnGUSudf1mpDFmcZ7qTeNR
kaUbv85hPQlreOUN8uzF9t2Vl1uYPQ6OLLZX91S/8Gj4NrtDyG1Gavjs3uz9XQMRfn4gsjCWzH7v
UsBEioNwPN9I+/EJsHiOGKmRpf2DT8v8kly3yauSCATO23Q9rqKnBpH1JbG2DNNUKgQhH51QGI1/
uiiGFuajxnqQrI7u882J5Q1EwitFGroQzGelFw0klA9sNE7N2RoB3qJdH9Wmcc3FKFw1Oh6m1723
Zh9sYYdRwwbvIQB194cenEPHQ2wE2xSdyillG4VXOYulM2D4x2ZIiV4hF8aDLzqg1pKecUJej0Cd
YYY8IvPbWjUukvItWQ6GCUR/OkIkuQOOAWvZpgTp9mYNRjJmHHSMAP58sdyDvzXCnzPIHbnE32j/
NdxuKyMM6fbpbBlpi98tgI1OtRvjqmU2CqhbH3lTzsFk3QY0yzLDxVUjQwiGk63el0AdmnFmmlHX
swIEUwa6llaZN/hhcvUit6O+vn2iFvccNT0ykPMGbydHP/x8cGoQ3yc3GwJZuUDmuG9R59PBDej7
Vju3tXxRDoj83SRuHTFZjRcm4kmSc0sf/+K9MVoOaMEYzJuEQ5UBPsrfsJxO58boPypd2tHtYfAa
jG4eClLkk/KW0f9m/hwQIhcreap3GskgoUSRH6qJ4bZq1vaOk3fRciQfFZiCedLF8mYwYKUHKmLs
bqvxDFiBtWvZjUAPGpl8AIkBtLHssUrGuNpwzpG5piU19R61N5h6snql08cexC9lKJQDDQMSLHjX
CEyZBPUMNX+xPq3Gfu3NTLEIkPxkACRuN01vAzvJBkB5FpZKBYfhVS3M2p0uw0pjnUIviQoyvIHn
7epNlKUqMBBkkXDPyXadTkquVAfKRLQVybaGcSgDhMZF2fDOhbE0OjHDChj4o3wDUrrmGUak+TIq
SZAQPupaC0N765ub+4Ty+zXi47IQLvJamQyNBZKTeqT39hRj/Yrm1qWzgZQCW4r3qqKcQLZu0GId
2zQGoUWATgandLA46LXwvPgq+PCjDbbMymWzPER21EfZ5VRDHm+OS0S1daAFKStQs8+NziYbscdO
Rt/VIvsuO4pwu4zT6jVhJQ8P31L51RDjNdjRnoMizJp8Y2InzurOM/goUl6CItU2nH0DLjeKWf1G
j9y8A5mfTw3rqe8SMXz87DLUOEYrdpbDf0OxYgZAE96Onz4jRRXgQhv0dp1671EdofhdoZfQXRXR
rTrzbfY5mTgjz4eqmnZXCRwrz8AA9XFo7MkahIx8ncPSbXEdJl1cKbKxQFzIK3WNix3s+LLylqg5
Gr3zHZRSyoHFv9Jch7RdxOU4XVfwOxXtK7MfYsSw+i2Lo8MIp0AH5W5A83J78lUmZK1DQfGIK9tc
9AiRcdwb5DZ2szS1L2YaPEJxsJptC6AtIzg0ryj0rs+GLwY5pMJOmbgOG9JSO5rFFkgnK0FJtSrh
BSUcUGcdBiRoDnC5HMxfuzduxYzl5wJCgZE9rexgf0IknsbmCXc/ETY+NBPo54jgJT8vhJt3cl/+
ELd+f7l8WXIJXFIjcRJhKN0aWVWPRogP7oA1EVfFKW9fFFq1AymagdAMqG43f1DaiwCvAYDP1W7p
T3e0kTGn2t4JTyioazeZuBjbRTPd1S2SjUyaIHidcxkqbst3KS6UIJd331aUBUWv350zP9WpmxcQ
10cdIpgXe9o9A/PVn/d8mM9yr5w4gNU4ZWZDrliDU2EHtcR1N1p0QsFtikFy/9g1WCUSdCS+rAM8
K9ImgreQhgrxAGpy1KRw7IHKjXljBsDxhEnAejw4eWFa4nCEO0qFHITTSxe3d6G8/sVEFjMv/5By
gG2Mfne7U7pUrTy7IYRE8XC6UNnentmIcMGA+JAzakzFdbwZhdy8tL06cvzqgyyf4XyU9ahY2PfX
N9C04W3Z1G8Kj4/sGaOYFQUKLLh6SfSJ4VomSFpVoj3vjRFrFcsgQD92Gnwb27nnn5DkGdTCsbgE
0+yg/4YGIPQYqeSMuOtpw0PdPL6joW8e6pxAntWRDQ9UMTvCCGYrh7NFu8KhI2CWKD3HyJZqrjeQ
EbIwMS9SMO88CbaLhg4VHDoZzdnD0KpV3eYmSkGU7awsPab8Czb8WvX0bVXW25i5GkAoN6wI4wdW
CqlTrnbA1Ab4n+OxT9zOx3kkwHBpgYLx/aoV2W3lmyM1SoAWbdHbNgGQvh7IEG6dFE4pXJCFww9G
lP6Ap9CivyhledUeGnfFr3S4OJPDkifyt559HOnYKq6DkgJF0k8Ym07Y+Do630Z+pJsUYe0V03xJ
VskOCYkXCZzKWO6Kr4XknuvMzNvVYH0S5McUy39w/ceMlE9QXXlqxJD8MfiebKsvGn20gU0VtrKE
RA018L1hjzYvKC9qcdyfCMqRLe5dLUR8EwV1pWlJEYCXT5BuiHDge+BMfWEpzhU3EBxTRoRuRDuT
ehWbNFbu32FiUVVmgDACIag4IBFAILnvaY19vrjLSjCe1j+la/183BLu14yUqnTd+w/mbMdrAyTe
ogyoMZsom5EDd9jPahOUwHlKgMGPuqE/54n4hYAlWpjb32wZ/F574OJxdSxytn4ZvCRYLhrt5ba4
uXD8EorsfUHB2tfydpmgla67f/LW+Ng7vAxRNpbMnWbsJ819Z09cAkvXYGO8QPM8xzZkpFmNCMOE
xqm04B5+uYPzt+PnQIOB53rnOdIHYgYvUtfb1sraHxARO7bg4XehlT3NIDrFPEGvfPDkgSjtwYRN
ilzRarJg5Kr5o5HE16/lXkoffSZ7PdyJS03eoQfaMnOMStcQ/oVkf4+FH1dvjgSMQSaWLBAJYOpa
yGIkOq5HbJw5pj9JMJvL5K0nDleEKF+rV+P8sVBwRAI/pyWQxekBimo8+PersI/ruP1+Ep+f24bR
hFiV1sAwIlKp59MP6d9SRtIY4gs/+DW/hKJdT1lTRX6nDFxRzvMdNZRUzzmgkPNesep9T4rK3Gmy
+G/uSmUKVGMsG3/unYS0ERrK5ggC7LA+keNLMpJ74dfRqUZIFodi0EIExhtaDXPLpSnHJnN6PXT5
/qGeP/7qXo3zxDx4MvSZAtwryW93q1dGZg7sAgU35eYAKKFbq6NEqz7ULjciGL8fMhKnrz5oL2sj
7ZttSa0EtvZqkKgky5bnTKntshzByJr6YxCg+RvpywCHxVSc+fWGLl4jQHnsiIR6AEm2NbA2ZiuF
oQY+z0Ts9gpeCp2631UEYPSlYRlVBdrrjuFDfdGwo3KRNz6H9DFNDOA+WmiJPG47VAXr8Uu8qlXW
AW6b573jnUY+cWm75MOtLvE8dtbmO/Cxd7Lrd4eevHkuFwctonlJeUJlmgW8cdXWUuIqigjJIzOm
DK8C1wMCXTu2HSWjV4TbQZ/VVhbMK+DV64puFF9RvtPap6nsGHjfWXgQ7taes1A1Wjt4rClX9yiq
ehaIARxcosR+lKPgCo3xMzmvET4PjNhUImemy6qHbtQxkT5b7bOoI/1cz6z1snWFmyK05zww49bh
R64kOBbT8ileNE1CizW3naqjwkwxPSk4k02KjcnzcyrDWYJTFjxNpN2P7N4QthdVqpFlIZ0LPlAH
4w+uNVuyJCk+lvFpalqx/OSbsJffBGiq6hPd0x6FaeZNbS3KMxqbBxEOYZyz8wMuuRK7ggT+GsNp
eSnTR670rXy7wUsHWI+OeQkro5S+iNbM4dlDyXzpV7W4k/ms7ykAEWz0l0MESXtRUPb80zSLLtPM
d5wGrAN0sf8pKjS2MnCUSq8H30Io+V8j8OgL8+/oaWAFjVTedEDRb4kcUWZaPYgwtKRvihvzZ6QR
9RP+VE81qVOHfdknA9DNFYVk5/jhcYGziyer+uLc12tFqIy4GCJtDeUMnTa+/DOvMwu/73X93IhL
Vbs/9zf5HXom6NyfnPwctVaQHVt8YRazKjFQPKSkPwOQhAKakF5VWrsKO0ewqt3PHv+JkLwncvtM
zOcVNazgntceJhraw82Wf7aatBdN1cRcjyMd2baveeP81jl4d0m6k1AvZwRGVu6HONm1vwxt7M/B
UaSncCUZAFeVmy6rHrlW6dL4u6UtFxV2hywRfKvmxDOVorUgARvB+ebGV9yf5051sb/W5HC2RYT/
HgJrwabuMjyqROs/O2Y8/ri5Uiz992MmX/YcY+xX3nXfQl2e2tAW0NQFwHQyH6eqw5ikg4sO/BZ3
CHRyi26JQNE47ymb50lQBhhEDLl6NKm1ugEQL2ewARac4U6y3FyTP+YF3I2ntxsXXysMD0MblR6A
h6AfilYEP4pWS/HGe1hXZclOmJOo5455Wc1nhdKml9IXPYixPr4BIPr9oL6O7L5qYW5/1ZD8AMjI
q76CI8WVLDlzhkIKKoxY43zqI9lqDLVvtn0E/qSgg5tBcfwOZM0SDm3krUNrGll/3gCqMR/Qc8EK
lAXl0s4XDl7pJ6xqE1B+TfaAVe4cb9gjlDoBBG7rK4FLuuxEiuJJd/U0zv70QWmHwPRSNc03LAiL
mJxzx9CqPecQOZxZnMKbKYoGzMo47iIsvkYWFnvkbNevoHsLSo4nhHV8mxBFxJQK+W5yBoA9VWio
2nIFbW+1cAD3AB0G6cQhNY4K15d4d6wE9xCY9+KuDd5vuo0XOIozy+w/VQn2bZA+6PMeVG5CvSTQ
6VZkjBcTz3eVLdBisulX1r7WxF3WrQo9Rw0sjrmP/L5/rrsKPcshDIWmDypw9MkhNZx4ayIAjHov
xtSCS3sT1S1zKthwHncy658CNUnsdAAUXUewEr2ciHvmBVNnVnBBfbgnA9HuUN2hhz5hWYCsDujA
N9JDdF5fMApxZrr0nSS/8FZWtxeNgdCsSsNFBcRq+TQ8Nw/TPmQF+W/Wc2moHwnBgvhf5JAg+Jbd
FRn0TNJlnc1KYH5TcgXzAr7XoT2qiJBO1pbO9FU+zFh9THG62oS+YU76NlrQHvUHS6sc5/cY1FAP
Vwgth33gLTOkv7fHPMe9ctWvV5NPrjq64p01gsxij/ebEt+d8YeCQA7x6/+aH9wMLso5Ep3Vtqxz
6r/ya9jfWtbnpvP/gJdnuEqHoJ3V/YswhtAYe+A1RpYR/X3834Vsk45loHUi4vnLsJ4QDMqAQn1M
U5tCj68mUJbrWgoaMZSxlw0BtxT9To92e/ZtmlMidFzxPM7LGA8jEOBIbUm8Z46+HKXoueqL+S4N
xpn/cWwzifsEKCv8V3SvAv9RStc9yXlHaurQ+bayBV4bryMow0vdglfnCh1DKtIG6GURiWQv4udv
WN/IpKoeyTFAvxWWy/cSgP+3xFLRXiFDat71bHID8ineXmAJ2Zc25L4zGSAJ6PFl/X8uyEn1aFmU
QeMbziuRu+NsGnI+M1i1ra49D1+6nbN6JBTqXab/b/ADrCep7vL+hEw2aerfUA1ccCsxNn5CYT9o
mf57NJ4jcjEJlkXrjJwyI0jsP5IlKc+GXi4HXjwuh1zWVpdZ/FVzf96t3yVhI6QYSEKDIQQRC17e
nk4U3et/te53SEA+Z4i4ZckVAf09r+gC9VBZPxGe/DLdLSt3TMRgOqg7G4KqRVq8z4AnIaH+BtE6
sesIhqyYoNb1qG/6JgFNXr3/jWulRrUL1MHU2u2iX6Xyah74w6lVqONzOQjHMg9x+gx7doyGcIa4
YcciwiAgsaZTdD6NoWQllhHmhD63FL3nAFdn4suJ2Op0pY7z1NWslGuM1k9VYfmPtdcC6r1LtUa7
+fWyGCCI6aW1Fk6VPlyA/1sfZNzGwtCGWTwwQJ7fPy18oYszi8BuxO0YPkc0qfv1KpwSmYO5zzYn
dhhs3ml1SEbvAqct7nZTL/m9t2Xe6I1bDtDtc+XofaMOhGlLZsxUB3QWDQmlPmV3Xn0JQqgBjk2J
YS0fNIlU9NW7Do0ACmUgZE5A9ZM/5zmRQmi6uGeasb6UAtlmwdRZqhy9yDVbcS5MZdbirm5n3Ljz
QiAyYS9rqV4e/f0XbUXJWVlKN2U7sjFPa6qTnD5CooZjTPyZY3gn2l+oLCzRbsWkNrFXYaVX98W8
9coo5hzvO3yPOs7cTlD1RoCiq/tUpUsA58Mvpp/9CGcfPfKJ9P1+C1izzOzLEZiDhS1KFWdlXp+7
oVDYUpwUBrvxq2oZ8oqWij6xnvQUYeHKHtYjNyu5u8OSv4llOS7lDbZtThDJsOFgU6KIesdEWAic
Ka5SBYpRBQppeY4HbxqN403QEE+NdyHOcTMLNqKoYW9427i3EkXMIPUlxK1NwEJ7SkF293biCkg3
pFCQHHPg2ojwzBr1SAgJSqtuThcXx2RlUGu6UX95wBx7Fjr5D+oZBMcPTDCisWhsj4whK0DObFNF
ImUjFn/z+5uB8UV1zsOkfHCFZVPjjdOJGqnnCDCUJmUJMPD+0M11naL6cYPdOVfpS2U9UrNKby38
RFLLnTV/+w/oSNw4el+hG8bwGKUkIJPdLh6eHfy1AqJxcrcUWKEqrTFSMaqmQIqY8rgDO63Q9xgi
/wU9DWOodvkznZvjRvx/BUOnn/KlPMfZfsXp4eo79PUDCW9Mjgx+BKZlV5Gmt8Lfts643cKpbEHP
mVp3s/pUxIWDNKMpTF1KGcDd08Dy6JgNamQn+iTM5adn8d+UHsg2Pey4oqh9cAn6pqVrSZoqj5En
E3RXn8/6kE/5VIy2lgru9Q1+ioCCSGDPS6ENcGEYYg4Q9s7lbNR5DOkai0g0OKkKzgGIGcr1NI4I
lv6PUFkOrjT8kpB529he9qGZ5yQK+IKJpOnhPAzubWt2i3JhicGaex19zMctj/6hmACXD5bCt7Tw
yL3WDV32Jbhq8p5v840oMT4V3xYbFkg+zg+G83WfMynbYGU19/iiIyNEpgEdCKuquTh0j3H1HSRK
dDfsofYm2rd2mCJyQMvKAFwU3lgqvXXlIT8htzJObZb/Ss15gw73F9QnVk8h/lGCM3saHNb4k0Gk
yzsgT38UmhD9uilOtgXTBpWfiKBEaLD4dqdQgSGYjJEIQNbjo9vqfq17GR6cm7s6mZ3lmCpW3drx
5YYOUAKqYmuh+iDz2oIpxMK+k65ZReBzahOW1CENQQn5Ze2L10Qv4AvWzpLIHo7FM2U+GuKzrFl9
bn6G7kxilJ1tR2h911hi7jge9oKK44D8kA9cZH/2jLqP6jO7N8stLPBjvRKtnwkzpfRlgUYEvaOT
f7hr3gZm2FyedfMMRnzw7lJJ03E/bICB/kTzOEIiihfEhzlTHDmhBL8e0bOtLzIwjetLU2WPPTT/
57b8NmR0Mxy3QnLirKqXPqmRr0GrQ/TIO/O/qESeQ4UBkqKSRihfnno82HIru93rXyANMRC4ACLP
LZVfnsX54/3BND7vSQQX5PgN7bGrbz5L5dmC98Di6Q54BCiphMSx+AwM3o8ghCwS7AbdtQ2zhi4W
fvuIBnPHRXyY6i+1+NQCN3zZrXnVJk2fjQaNqbSjbsVzxA9/vf7cbYBWQQRh7II+05dMj6D5cY31
JXWtJJFBA2rOzoc6HwR2XbZhZ1jyL1L7OAqVB40opnma8EJkun7HWEoy5ctyGZx+fLNkh3ys+5fu
4c9qa4mC6FrTq7JA+8gUYjiO2om6Gj9IiW+hvZUqIUdJfObQ7XRTHquYudrWIJUPe/g0uSGRSEeC
EDHkiBqiYfn8eJ/yU/CVc2471QIZuuZieSRSsQpl/GCVumrda+JB75gCJNURMD8Q0h0obwgqub76
8NKecsG8K2WB3341dS+tjJsy5G6GZ3heHZ3ijjBMXBehpqlsRm5Gd26YgUWJKoGAj6cfekx69W/J
g9HSTwhuEXwDAoKLlYbD8ED6VRQAAP4AlwYc5DCz94JZxmt8C+ghwpKkx/vOdLqTzFFqaA6EUKGd
VQUG+7Rxrw9XZmPXZaKz3OPSae1jaU0sKee3aslB9pOTjm8UwJT69TP2C15/1SQ+43xkSb4YLplv
raw/UZiz428wr2tUfOF7SoZwX9ZXGwMVNRbORQi4YxKKcdP0euUdCCIkdjuhbMc45F2izuBGBzCo
CSYrYPg5ZdtcCoAPue6eMhh1JGyP5vsxVqcXp8sfQfYqhwh5M692m6OiQnZNKwyyxCpAsH0SNx22
J5VBI7uu29C4q1CHasO+U4YeoJCXU60Jgjvn8ynmPJPi/mC0kICvJEiBH+3k8ckoEmbpNysBvlDK
OvzJPkW819ZryLw46titYTzWWvVN/rocWYt/hzKnf8g0IJmk5YSmiKbqT9XKrQU+estrTHzLkpXq
5lqvaCGgDzcjwZjQ473wMdOdXGMIBaoZ7ZvzJd6sotNUZ6Kap9ZT8oe2tT2uuhZnHsrVGgZWUCak
EBFnhVzo6vylq5yzX6dzFOFNYqDhpdNT6DpvNx8ffmaLBDpYYqmaSSaNqFPrhZJ7evaTER+51lH/
WckGOIhiX7o+rXebqiVzLS95FhDgYvYjqhq9aNRRPeJ13Ws9IqDC2gj6b9Fr7e599QBqF4pxwp+t
1/0nbspNqiM/Putj69pvTIkCy0nQE3YuzdpOLeiAB7vSr/af8CuP737u9Baes/G76RQNjNxoSO2L
qcV4FXIOHORkAqj0m20tA19MMW/M+/CZxE8EaYqh0yJZLyL71goinvuBAAWuLhXHN4oYgwxXu6ie
TAxk+PdC2U8CxOYEXWd5EnW/e1AA/Ol6Hi9fRPAggwm5K/cKleq8sahzkgAhul4b2WP2nKms3cbf
homOwuu4gKZYt1T4KeaP370zmhet+PguzbvGnPjl1vnSBKLA3TckCOWUQUqKMyF2KkJ7Q22+RqYy
qUaRwHEuD4PvnT68ROqMOewChTK5iggxga1bE5vXtkkaZIPDabdv3lTsmdWphPxVGdoP0jY5Po3S
zirqVWTcLCjOu+bKQAWT8BKtqdm+tjMdUGxovkQy7HKnDyoZ6Pcpw80Xt4TT8Ux2NcB5AWbo+u5G
QpL3gpO8nWCOEk++s0KeHADGcGavCuxb/VKCjVOp9dJ0yW8qLZRexMlVpSt5H0m1R6wyT2ur7MHi
JGlUGpXHbnJGe+bqehscpaLUBAJCxsVzdvuhPvwD5Wdd3N4FCniTbh5JMKO9Y1FG5y/aGegudwkc
VurZyOh5N8Ss8jm7rd+RVEim2yyXGbEbUET6fGlATuis6fA6mWAx+TsuGHKX3pK308ZkbUYnwO8u
MCvqJBqRYPR98cxzleT4d8FB/WocieN7vtbzlip50lNnkpXIJHNZUe7VfRxF+CO8XinYkihSdzYX
1jMxNiMjAvckpkjpRjCQDyiFt/nbo25bYJzYjE0AgsMeVjk7GWoRfLMRClSFzWzX3W8xYLRvUeLA
3ZnOg9rzRlZbd52RNsgjO6bFhn1wuBwARupsyO2qOyKnk5EZ+r2m0FVm+qGk5fv+8Somudf0ZO0O
Pk6+mbAekZNiGgYqCsPdoT1FLSsY3numYrE9KLCLADwjEtMEXPV3wYiMX+sthWFn2uCKYPSSaj3J
P06qAWquAKeyE0hAacdWDzeDL9VxH7HWQMhu9QqkKIDewjiAUbf49WyEuYlgZ2B3iznQbR+zhOyh
2FHohrcPV/Buqu2qq7ZYmh8lLge9H972pmx0+vsDrg5uY4TtQnr5QBYyuCULml3TZFVeIlW/yI6c
XcowyTBjJNwurydyF6R0ONEJPYSDYY33Pft0PPOkRipbBqTUwmTSEAKUZBl/X42aLs6sPwNdCLqp
Xw2i3xCTW5igneLInG6VL3T1sB5VR2krgolHkgBBwNp0O/aqY6uFEIQ180bgWTutydGMQuMBWQ3y
v0cmvLHBBel6B1NiVoCFHbnncNjrdYlSDceZkOSAqltUxI5OyWzIm2pAEVvH/EBsJuWXhwKf8zGu
k0ZZu/p7sZ5CmHcdanvL0JI7gZvyEo9rBs8fCvseRuao48NCJG8DIa3HCF538ypIqiSgkQCa4/7v
EVuTmNH0V0cT0PMWVG2RldrgyIZx521Kn98/JF8TZxAODsngpMQXU3MFYsTENd4O3zrkI0iBMWK0
of8JqHw+m/fzzfcb1ZRCfKrQAXwQ4N+vn1nGujbNoMt90EAvRVl5Xw+vM2cG/LjT+mTvjZeb3i28
rkAEiG/f17n7KBlklzZ+um+o9RlJ+AXREfDQ/yJ2pK6n8yYW+zATwh8qeBdfAmtYDNplSht0DV2W
cNfsYOxRBL0ojhoNuO1UdPH8bw7KHfAdMvV1tiJZLuHyTZo+gQTbTmBTonbRL92kZkFwTEqc+sVO
YWzlmevwm8IRBP2tdaR1pOs5ehmhB6seOSixpn/vE/WjUsZpPxeZhq/f6iSw5n2frvKcODB4cVLl
gfkEp7iPdSjgAVmqhsfz0Zo3sv1GjvB2j+J02HPxAQfzObgFfnr9RFZ6VsRAn3XfTMLV7KBAwC2H
Fj6UUmm29GcJ+SYreLc12AK76wGta42/pS5BnshjcGu+hK1UmJVMHbeF6GETLRP3lmC05Hdizfh3
yvDhHVdveXhvQ2NLB15FdFOOQTWrqcRf8LizD9Riu9h9RYaGSyxMZZwC3MTbFfcNE9dqkHQotxSW
XQTXVxhLhrGsVVXUaqJq0tB71S0Kb+OclpVsUQFvlB3ZBZsLPGjX2Ercd4WINwgVj63hBMx35hQC
2ojM/1izfwPSzGEZJc3VxH9tjaEzy9nI8WOPjGODeCwor9XfKdGzByZho09uQnAqFLDvQyxDKo02
H4te6jgKc30xjk0lBO+84XA/gQKsfmkcHh/pvN3Jn7qZCZUjadwV5JaOFYsSuU8zcCRqS1YHJUOe
gM0Ek3HuwtozRbxYPhDca5YZAbOZ1ZI3UTNrmTJ6oMn/EGPBfeYgh8sCGACOynZtG6nt43VITg3Z
CkgPHgs7vZlwyrUotNtj0I7OLsv19zFNhUerRp1qetZiwEwPnrxHHjQa6Itue01ecHLe8Ruz5Ieu
goJOS+Lgi8P8id23FHY38nneHk7DA9Dlp6mw97SexiV6FxDFa9nxc9n5/iqb07n/Qmjm40/YXd6z
U507ZX9DAHy5dQHpHyXptsWzcxbqbUM4nwoGFXbpglxfsGkc2ZK1Ca0IWFRnzg8putBnqnC5Ct6z
dZxA62bTejRTJ1QxPc/2KvBqzhYXTXP+UdWro6INuCaHlFYfG1Qmuk2c+VrcVf+bLmHpfpJPw5AK
4U1sZRJYyE7QSmf31UdNbXbq/phyKSnIMrJBbkS3pR9pJAh6uYm6la+96x+ZXOGG2k7rndlJDrbW
StQZ51fL/jqDNBG0+2H0R9xYrwD4ywmyAS8weAIXQKF9ITGhmu9MeqC7GfaXmU+rbPR6ycnYqqNp
xALErQZUuAxSTo1QgBH/xM6ay89kJYqkLt1CnmZy4Fjhs43aMgiMFws5yX7jtRm4Ax+MtsViq9b0
RQjSmmF6kTxdwXpk1ggY4IKwptiC9USAGCUdDCwwdREJfIS8OC2EZ8xmzOnC6EaiMRuknuyX+McP
kw10HBa1GkJvyQwfmzth6mCx+FDgay6FcstwIMesTO07bK9rKK/tjY2FvuMp3FInWlCP2ehwQF2I
Z+saxlklCyRY2dZlBg76bMAT6C1gMBjIq50hX5xufXqS34yGv+pD4yBZN6hWyzNhF+S4tTY+Q2Mk
EfS7eSdHNdR11I7YKSRuBm1rUMfoVbsrp9sg8nu6yv+b3tY6yHHGsTa5oUhPoRe3P4PGR8MyXgnx
ZD6QkMkVl1yJywlxVENMbQgACM/tkT3ARsSVql9qVwObS7Nmqbb6T5a1n28eLoyiZCYOBM4VfNDb
829DRZ1D0V5mb0WMRZJbDVwJSq5EjGIt44qiEMZ0gQ6fMnqviV2mB9BNE0rz3Tt8NB+n3joGW6bn
adIyE4PSrHNivvufPiUMtJCxIMwXUBRcnOC+tr3iKAreQBzx1iZ8geja7GQ3IJG5t1LLIulRnrBK
avhzGuxh4eSw8I2xl7SFzWmg0WBpBXptORc+PQKgSyyjG5ZiVZuRm85ym6R1Ebey2PcfD2J858rp
fmus4OdnfrXM4/JtnHq4+O/U6tyFK1BIdvLfFDDR2woxIzixXyL6dLZGlyB9Dgzow7x3JZK1z4Nd
wrwajIJ88avjEEjWYGIpP8zEyfcCQWLrEx/15c9DpHXZmsv5tFuReoK17bQRXXSF+37qUyprVZB/
fjlrTtVUnT1GkM+wcQqsAvCmTbzpUIb3qGtjNVda2LAvXIHTHWpBkJEQwiCfnVP4X4XQwu1iqana
1VO3S/FtsG4haagLkbEHmUpc2f0mhaffRyV1z1TFMkweagCi9Bludvhw79vH67C3nm5gK19IDqOc
7uUQhyIw7QJodB0Y4HMQwegoPaV7JK9uq9qv0k0TnzJY0vN+zH+jWxnBe8E12rm8EK5uI8jr2F8y
pZXLsvywYdR097L9y7Onz0X0TlTGz1eititQEi/UrF+zrhkQ3J1E6fB/+pcOqKBpWe1y/gl4yzgc
SjCOA9opCVCeIKQpU2vn5B6ExB6SvbFWAOJ8dNkOZA5hYOjyFpDvQNG6J6YT/RWj5QuxG3+2k5h1
TDiFFdRkKVibpqX4V0dlpBl9pibsQJEpe/7nH4tzU26ZQJH3AYr20mHCpDa01r+/g5cngq76FV0j
tTYw+HaL0623dpxu50gB2my1R3nGbAWpQfvBta2hIYlQ/ATMvyWVZFwPKYWrdHcOSaHXwmZ2gOuO
XBiXh4USt+0uGZbfc2oBSo0xWkH5KC35fnpr5wsl6AeYEckLqtTTY+JocaH8UWzCRK+hmwX5c3Vj
aMRQIXD/DpEQH5ptb540tijTmhNalchsc+2JMDbFBGgXf1eHyCk1WtdRflzzrCV37oVDexFFTGlS
G7BLwcC7k8KdJxzAKboW6YAk0m7EPZAiPmQPW5OO4Ts19cD1BFNPIg0hHKlVcmtnXl8zh6T/et+r
BFqhC0JLlsCmeSgS36T2ipbc+zDttdlCgVR5Rpm63c20HBQ76v7DMuTRsn0ZgOlgEy7BCTvJKd5V
cvAzeqvp3fa7v7ACi5K5zVfXwgF2lZNKaKwbcRbzVh9g/umhWjqPRzUYDprfRbmD+3RAxSpud+mf
dud4PfFR5FRkSOUKc0VUFPFHxlsAj+jtwWH1JjlpKARdDtNeuhoun94PZ+eIcMp5IpVY32llh/t7
tnWoPpSEai999H1dc6DaQxLRix7I+J7SrM8XimE/UHOClako4mWRE4C1Y752RAuJQHz1kdr+2sZy
DURk9HLHLySbUaB+Oj4YC4K1lehTuVzX9HL9fFmmrHFqOMu9j9CmX3ZU+S6bQfTZwjmkxzvLLmz3
HB20zv1q0FyHdVJHeixo3LskLLmiatAQT6cBIWBt7ELRoPi/+pYrrhNH1zK0GaWOmVRHOQ5MZRLW
TmvVBX3cN1VCuT5SEiilZOpiu9B68Wav7NqjtTetvXEmtQnzDiKlHlwlwXT5g/+i08Yv3P8BVWCk
Ws/gFrunXih2ErPGBFB56EtHIt81L1bSlEBTrTspWVrspARh0yR9iPbNnySCFT0Pgw1/4my2yhYF
E56KUDWrY5B3ISS5v/w6bcSqOmoIcqMlKhkkcok+zHqXvHE0kk5iATKKR1UMmiNWb6Uwgblsaz1Z
mVmThYvcGdObVz6g6krL0npKQVQO7PCB4Krmp+gc/lqNvf2tiwr1ehmKjDkbgU/NnacArZNnhUKi
dhXD8U9Bc+lpLl9Ki6Hot8AkBbe5PCoya11Ak10/BJzVOyGhJQNqK03f5Pn/ehyf6OqOZSMtUDr2
RH6/8rnb4G5GBOSqG+obxR84ifTY/mxnvbXZqPuJFm9Rnksta8yHgMtAzTODi20nnERYCNwEoW9z
hFo24bGt2qAtS742F1SnZZsntfijoe0aD7tKraWP/qK8276+IoxBZVe3MCEOcaNUBIgHEPd2WsHx
jeteIQIx/64iB3Dp4e3qTdiHxi/Zret8NHn/bQjNsmkw52opkC2+wzsV+5HAUdKGKMJfk9sQ13uP
AQryn9g4M/gV2ygYmmAyeWyOC71UoEZFumcmvwVO7CeF9PEuwrNKGxJmoKEMCoczKF51tBJVEqYk
v0a3ay26+L+++mNllhaTdSf4i/iTfyi+EmIc/vZLiJj8kMDamSFGWWwWqJZ1WC0dhkq0czU5Alia
bJ11B2no3/SwZqUYv9gE1WKuhRS8ScNpLPzIkMYyeRtC1xu4bDTkcwPBk91qOh1d0W4s3hHnaiwy
EHRs9XU6Q1ifvacEqzPH1OqiKNevTkti1Nwutmh+a9hh999Uq4j85IjcwbVIzEXcy2H1XL8QT/aO
RIPQQ3ka9Kj3ATfLehSIbz8lJ1fLwE50ZUjDJK/N7xbL0Bx80m8khJRCg8WlWD7vx8+9ObGG0Qo0
qQHz2tK8svNSJIdGn7GtOxuatxhuAGDPDB6BiQunabYqmek3u601WzDA2ipyV+Gtp/f410Xt8ZCi
9Sw/10InZEuWfDX5PsPU8zuYB5oCW9YYbf3SZopL4pMeY836Ikv/OJV5O+Yjv1P83DMc4SKt7yQB
iy7GLZaEBVwoAo2ZO9njHDHTVTduFlCukld0qsAxv3nssS/t0jrc/BWEw4IBwf8VEBjUh1au4Cej
6CAi8QkyCC+gR0rojopf8/yKt+oQ6nbjhr569gABJnwOC9wnJc37BKiOgIKMD5dwPjlmmR4e/2wO
JCRdS6tTTxf76nmKDMNyBgx48B46VBETikLhy158o/lQF/FLVz/x7KEuFi9BinYWf2ZM2dQK3IJo
nTv2K1hYraLteu8WVlLHoesQJj8iF3V8yXy/4N9dQMKjQL8eW4o8wKLafCFMbCYAsX2fgTLJ+yOn
0tkV79gAteiPWrfCTZA5Fl8PGAJoZmUZ1W1Y4CnxIS+5PD42nvhkvbxElvmr5pi5ORsZKBJ3GghT
07ibiXsQb3aBYt9m0hP7n7QByzY5Izssvc/thI2+6HDsadbgmVsw4jExBtge7e31UmAOATI0nnmH
IOdEAuCQAOlzpACWscUkygVO/1M6uk1+/sR8jD7YP41qd9ah8HLgIC/7h592ZQO+vx1lG2rrrD7k
OGzknSqljqUQ5t/RlW9nKnHaAN6pdWC570gBnKvmz+VCkhWAKACNN8KlKzW1+qqOT5eJswBeRllb
rM41gSTQ+f6Ir8VJQ1lduRss+Wc1zF4ajnxeLlQH3kmUfMSO0SNHYy0wqsDrwErJZWJdTNTioPpN
qhMhFY4jBh78BDlEMznCCxVyXSAPVQwFrT6uyHTAcsX1p4dKL+s29AxT2457NIzG2Dy8vAYSVk35
cVHLp4pTauBCjXGhgUW5KsEtNIbm2z/4e7Q+A7r+HNZMq8/DDjNq6zHSldE3vcx9m8GMj1bcyjZ1
8u1rZIuFSXySBZr/qGI3iTtw315Eo7qTYumexHMNRZevvefsDDsgg43KNjBiL2tia3b/hmrUWAo1
JkmhlivuCASaBwKppovXLxYYawPwGS/2vFxdnUB6I1VBmladW4nDZrmIHzAryreIw+JF4Mg2w7OV
/bWyaWrE/647IKzbqwn3IomNjmptZoCt8Qt4OzBRMftMemG1MATKldiP04YySxaZUPpcGVjzfip/
SEjWC2G9WuW/NHCRCM4/IDEoKWIMv1hegm9XsDD39GJXxNlkG7BOnxxJZKBaHCMncqsZLVxud1f3
pKG4Bk8xcJywF7TPB9sEVuucECdg2DEbHsTIb8XdkNUXNLVnfK9rIHalRKnHq1hg8Cum+qdQWwDz
nMwAJklbPfUKaEyfHvOqoaai1/DIUpc4oih8rcT6yO+wpEFKtJt9J0CcfSQwb84xJSlsgkIbqHcM
ktM/UhSmWd4dSn4OZsgOJfDOOzvmDB2b4yr2eghn2BDGIMPfU+WxWf4shZd4AAVwvL5aPDdjBugr
TunfY4NWfy1DyiJkamWkjkudmHkAVdwEy5ktosV73HItyDxQ57a/F5NVfMxHyZ99KJQFtsGcSSSU
YvLfDiEAK6Y2lCPA7vfVbha3CekAnyhHOp1gYYVH+dUqjSijxoUxa4OmjZSxS31pgXqNqlepOPmg
WzgwdH9Hv97mr52V/IiTYdXimhVtO7s9a9Ij6jV6ME2xtr37rFSEFWRqUA/CD7hfc9HAyiSI3pnG
Q36VE3CXyij2dwbcgZ//L23WVKDeaDfGj8rGJoGZk53z8VyF8wMkYhci9E2jc+VGgRrktyeNYo1L
GJB6GbQX6KR+YhzLNTwp0JQgMZPn/iDQSMoOccfUdvRdvMP5wBlb9fyQbBF7UZDj4fF2unHs43rZ
Rvnq6tcfkETcNynGfg2AdgUq9jLkpOGZZmBln8R3hqwqiJwD+cdiLNf/6ilibiHFeac65Atc9hy5
UWUjxtnENblXSkFCBnHiMR1jDrUUioOTMN9x76G9uSvresKJ8HmLhffjUqEHcPkaYRL9qUL0Lsmj
T1IWN2orY/deqARqUmAy0XOU9gCbLlWFXroJ9T27jfAiPJOo43J07CHCfJebxeXJyQ0xdEwT7bHZ
S40EnhkZW1dC+P3uHAKZpFPsgBgrnrWqFa0m+EEGDo1mibaq9hQHAALdW0HmBWGmSE8NzP5NPcFP
NOhe7cSbKv8ogVEUjT8cviUib9HIe/MbYJCo8FgOwwaUKvsohkE2kBnIaYJr3WNooMlCGVnJZmfb
YYHLql2JQfB0UFOemrl/Jt1WX/cWLnTRt/D34PMce7SIIBEcc7EOiOewXQLSyBcEI9XtvdJMX7KO
wNuFtV0Tt4oViyaFW8FvGTRkn3ngkiJE1r9W0duBwnSSy/Hfj4fIFjer4vsRJZxFneAgao/QhrL/
+XSNqkPY+5tYbGk7T0UXyLVwPxNZwTKD6rdyUujn5cZ12zn14WzkeDqZZCHj3vKahDQp6qhil6f8
gorfqDy3fyR4L58H+wa81Sx++EolOlcoaXtBmWz3mL1NFjU2QYo4EqkBT2lOXsuUJJeO5+fZBPcZ
46rJ0VXNH7r6DMrJ7iiDfDYYNvPPS+3f3df6yUeKa2vghDh3WUQg6Qlh/+GXXGdMXjl7yAaoev4e
OsSG6qMFJb8AsG85BlkVo96s5ugDFsZEeCAxhhYH5YkfuYIKq8+8t4DzamcB96b68s4v8Y3fwCMM
vpt0xgXmgNktlHCVd0O+X65BLaFW3rb+nGg4P5XbTmrh9+cn8osutq/v5mcaV5R8ig/Y88HhVCfm
JsdegKCnITw+REPLT5+ZiDJ0mL7+TsvnlRWv/9y9yRMvnUeiZB3fr/LkRz/Aws/gICUmqVtqlhCW
q3XUbXxafO+7at9eOO7yb0k3c2qzYI6Dk76vE2f4SeLHgXCL+iawyNmxi+2kDoRA5V3sMyW3K5RQ
KqvN0MuE+cxs7rOGhLVytR0e2pWwfU+bqVSIjkYGs/lkcV7eqTYCuGSB0D4Ao0eGq1ih/dsrbiSH
5aDj3e3h/q50gSvUY/uSc1RUTtLE9djajoLtjpd6o8zPSgedas+foogZPYm/BalbyfqLWalWIQxW
17YxBSWUT5oLeH3edQQD4FhVnNelYn68sy4A4ioLoRQVbxWXAsXejUMf62Fh0LQCLJ1Ijvlql+S/
P5rcJSogG804M2SdIInDl4EzQ0WRsW1HbsJwf3kWYXSLuOez3FYrnlGrP34IBiXd9cspEekBLgdy
CePeYwnb6DFZMAcHFhg8grTSelY34FKOWuyA0hQKmiDTx7BRjlVrKF6MWz9CjHSSwMi7vW5F/qiC
LUeUKWGeZSAY1OHZOZ9g7vWFB/NOAdPa4PtWNalvrZI/aQE8U1pQ1PaHJpZA8350IcR/O6Nc7DSO
MJNprFpj3J5SewldDU3aG42fWBM3mve6xSl4IcvlIob0jc5FXXQmjoUDYmdTcBW2E6jM3dHPyr3W
b29YTZJnXVyHnHxe1qBgH5dko1IqTpO1elgb2EGTBEIZr1phJd+NKUCxEjooALGe25EyIALECYJU
14lS060dzjIQX5vqMIUbCRzaWGlpSbpqsNXwrUd7Hn7CQuz0cRfGC4yhMwAzlMbBzFAkn7daprjr
fwu7K40i1oOBbXVFgav1G5iNUDKtybV4mGHx7BYt7+ETGtxNNznzXSbc+JskhdTyB5mgvJxFKVu0
KzHNU6T8dvJFyl9WVmWz2PZQSGY0eIDn79j99sPl65kNJRvnvEXAfx2651u8ioNWld+ljxqyMd4a
/b0Kd31gGby64OkTjBQaBkBb1l6JJKjNjpG2HJQq9Rz0IYorxXwF7YIp+UN3fxkn5nIsJRTSB6/Q
BkxFoJT5ZhsjA/CWT5zhFelG9RPnpNt4TTh9FY4nlHSO6E5ty5WLsxWXXUebvjseIpFvKlXLYnv3
GZ9XgNcR2EFYgoAlkvBUdkgbLAzU7DtfRUJ9yr7ekTJ8XEJ2o9nh0G/3Ltw+ahRoFvy9r7kAVebO
LF5a+M+cy3t8uihBgk6QsFzYya3HDJz+Efio2l0lhmMgiuRXv706r9xDFDS/DnIBg+UQuR9ZXjTR
J2d3EkJeoIPD2NQW41gTcjMhvnwNxwtRERlmQEfqkarzkU+FzKRHiV/4ln2DhBWqPoA0yeF2DX87
YuLmLcYXuy3d7VJMZHmxPWfExzMAVdrGnW5CqIn/cXpxc8ZNt6Dwjs5vc5rIbquWyyeK/ij4Azdd
aKzfYVDW40DdsKUFJLNhydyxPS+dhebxsJ319lhZp/tljIvKRfXnR+8gYQ6ib30f+s+vYhFp4Gv6
1fVL7vnzpRQZGygPA9eFvf8d+/VC9JeRtlP3gfNG8Kv0atR0+sn/Rl8MkQpmKsDFpEn/MGWCdYIA
OmRGpKKzuWJS3ebzA+3rMOlvkLrAneXe9OvncQNtAyyzndy4gZU2NTfJt+mCmVOnqgm6QuKr//M0
tD6CeCyVS57qDvFIBpGiZUxPDvqtO4a5XSDZjf0hEpp1plWVQdILh9YN527OLlWWNxw90ASReKez
fQ5/F0VmE73hNQOM5JrjzGv9hdPGa8vHDSUArq665KOlWIPqamylPj7tuf/MySbYKEf40reMrvsE
232VTzk2lRkOfOKKbBT6Ko34DUO2SbIjM9M6UgOInhIrggEjac/u6yNGiQLrkkjtMOoq736CcjCX
6mPf8ZzdT9ONRdl6kU/pKZy5orIHTZ+sEE5/xDuNJ2YcekJjMlpPUZrzWQAc3/mYHNusFG5cDb6M
ZNcruaB+sjCv0ckJEhixeZyetU3fqKd4t6CBTuvFizZQEDZ6OLue9q6++LzPVrq08kxFjnzhfIBN
PopFNt9Tq/yNleSyHIt0EO0U5D9mNL+FjJPP0Zwg+lOtaNJbRwjuQHTLWqZVBGG4JvpTgOvFNLem
innWg/svQdQYfbLKRXFg9FeXG/Q5b4e07oenqyj8U1Hx7QA/S/ZrxKYLUhR0LWUytuJf6WcLfPAp
HYSQqv1HdAdB78ZOs2ZiyJPPbeU1mp31vo5xxX7A2Q2wV7M2AnM0xngYJ3VoRDMiMf2Tm2zEbpxc
WVLygP77BRmC6up2VDwT5N9GlReVtrBco2ah1z4nbSa+hYsppy1PLIP8OPSzDgOhbzfyHaSr26WZ
Idc6qZdPiZSRTTCF8z13SOlQ8o4CaSmtSF7Dv9vDQQpusp9ryBML/YdU8/Xa3DxFTVKucX8KZdCG
+C41St9l9EuWHHLUgBAJ1ZsEQpaEcYzIGiwvrfTFEwQdheGGu3Q9Fl82lGf47fmIBMRW0P6GKjka
27vh4mJ//kNnECUY5Sevp7yMuEpy4rXVF/y0vCNTZ1ic/UOO4bYfGSI7+vY/J4lA7C68qYUySdgi
FWr3Trkaw/sfjJHziG3vKZYSqmTXIhCNaWGg/4bzcevnJLYEucUYU5AUJ43dRPDmC5LCP8wZyH3E
GZuLT/WWkVeTMCO5h4aqAXhXuiko8ooGeEr5WrNdUytzzWwHNyh3U0RA6bgxIR1obQXvMjQSkNqV
bU35OKIm8qTkAFSxwvf66Or/H4VfVaiwGE+MBnGpUcZReiFyqIHj5Yr5OPun1wc6AiWzr0WT1dop
TCqWzgS6CY1M+LpwwVZZc12+Xjz/BxqqjAYZ8OjKp+oTH/zNjn8wL/sSLZwkR3ZPtWwB3mO08rt5
Kn33ACfEz34jUJlfmRyfGBcIaY+/TDLbOydSKhKcl/iuLrRyLoI9dknNQBWvy8rIG5SLT5kzTKR8
/3JWeP1WjFEAzep/QTRkxaW28RHWwru0Xoae87MiCEzkVBW/kvRQZTXE75W/Kcp33neGHTKi5kNZ
tgYQk9dqs90dDmUAy3HvRoGdwEwIwwnyWgk3PEg1bMHFb2nB9/uuwz1IMUy+OOMmE6pBQxHbKf4w
i07t+o5ft5/Nahc3a6X/7PjsNQJ7QVHHgLMeyRetq8z2h8lp9fd1u1afB1dAdQz1hI/FKkewbgVE
UjzT13wuU6T1VOQ1Y5evc4sgC1bWleWF8BoJSFRzE6RooncZKurpojFTMu/w7huSENKzJTIi+sSL
9xS/zjrAe1l8TVLTBn8/u2nas8P3405ODurrpCzPNe3mwxiDdAqHBZWycYQfuuYEfvRlkoXUGh96
33LO2nKfLy5V/vQiOh6EeXfxiO96pyF9kRxEMT5JEVFW2HHBOQbnEJOdwQvWnSrThApPv3elckJz
KPFjHE+8vvqR5XSj6CEOBRzVR6F19Tes53JLm7CJNnHpAk3zkhLfRDjyaRqkOfLEIWxJvSvzugvO
vsdeaylsXCMPSXxqo12Sl2WQ4QZfB75tsaGBf7Vdv63XEmdwcovxnbGX3kN++XFUCOgcAxewOik8
KNB8Hxs6NKcipFPjfhZVE2iRRPL4LYG5L9JD0ObmosPDlKL69dVIhtnWhqSFMwOlbxhJBRqCZ1us
qhNvH4s2TYyUTeFdxsALe9zueCLVs8rBsa5gX7z/93O60cy9stwL1FJUcx5kN6H4RL5k732aYA2Z
O2PebwljgISPwXgLQNnQ2UGmlrxRsPcPt6Z2VS6/T7m9b3BYSwTzKTWXsYRVsWESy/Co4TWLmHuw
bh8xfwLr6B4g50YHBrd55DWL0OfGhIxAMhiJ/vbgsdxgMfHaoZFlNvE724x+zvQv9r6P5YUq0/PO
uOlB64Yzj2aQNk1hUUf5ISa3p2Os/IS+NsaNvk7UEiENFpme9ySMhkiYtyZM9miS4oxJKL6VXczs
9OYpFUok4Lgv+o/AY3lhDi58VYiwJgIfUmfuhesfxLRthq4Gu342RUfZAi6C9J/LP/9AgOB/ZY++
5rDZKm2GiOp5wbAeNCarh/JWaWB0vcBKZ024vx3XCeNIn/pXgBfLMWpSCgQdol56EJdKxWqEdigh
ZVdjiAKfqnD9ui0QMrGYryqro0bQ5sfilx+yFkPB5G3VAbNkyivZ6QHvh0rHEZM4CMmkBLSaX+E5
HZGM9Tqx8j/FMQ8Cnw9yrC7w6thvWoUFDNnep7wzwQ4cBmo0tTtB80GMtw4oe1cY6yvrD8fhwADu
qR0vqQ+7uT33BfwJAW9dojmxZnMgTEUJApDqZpXlp0ERbWkR6mUrQqH357xk0rznfxoQOGKGGzoK
1sXT0pLtsPOfNkvMSSqg7SCkq6f5Yirb+Vgt30ILgeuoU+GX0B4IrTPqZWOS1426vAfMMFBANP7N
8IBFCHlkIjVfZ7qFOupCoVW1uikOH0vvGqif4RqNVKnc6+URi60dMmcU2o6SYZJHWZ+CGLLT92to
+NQm7ZyxkQ8tWb5GarhW0h2QDCGx8vHdii7H52T4pUF59sFQN05NUoH622OKZ35bj1BWRjLr8ybf
FlUguB4HdT4aOorskYyjnxcoH/ool1N7FQQkA4sCml1eI+zWUz0VgOeHj8wuJaOZvlZPLCTGBijO
qghkpV+OUeY9jyr93+YHHOtlYZnrjlMe8wk/jN28e1v4Ni2QHbyigdSRIWNRglB8ucr10Jc7eD/w
RSYZgoYEt5I0SXIpun3UPK4yoxeu46d7ly1c9iFvKDdbkKGEzTm/oLSUCINOdvooc6YzK2vfElUi
//luvUu5vacczoeJoDgSPl7BXN5P0/juM/yRoXI52R5q9lMvpx67kNC0yd0hbUrDHIM/L3lZln+Q
gCOspqrW8ipth8eKdl61Y7FiE1UpFqWR2uLvcrq2Ho6jmmSKHroCdu2ROSf+sf+cY5BbNzprjQO5
1Bzvwn/tSi3UVLs0LljW/rm3ANRlKxgMRJKYs5yTSWtTr9gm+ugTHQyD2sWQWuHn8+O0oA+Tmcc8
t/8E23CnnXMMfIZoHovWdg64mzsIkOdRo2csdVepJmJTIfn7kwL1u4Cvr3wGvKMAaamZRNXXHwZ1
QHZbt95ZaEx5y0wdi4v6j2QLcSXVuI9IyD+NM6oiG4Cr2AqbVzNUTMhbFsb0ZODcDutGWDtIp0IB
9qYj2cJgoV92czTaM9tyUCKh/j8asjAP0gerxetfIbjIdrK8YyOBCy3rMuP3TmZSKJuByhJxsx75
I0LpmgWNMf4FivxPeZ79WaenFkT+z0O9joQUGWZVfy1PerzvXxXUPxC1mj1rk8sFVyB1g3myBFN3
NgXe4ionw0gZs8ceacwvnMlvZI51RMpT/50EM0VNdfiBqZxKfmLYdSn6Gd/TdoBDWXJtwDenLXR7
g/8RXQXoHT7hp2z/+h3bsYHaugkrcNTbe7LaMc9ZxAtVGN5brP3/QY2RyrCv+leuCUXSRXl7xNFu
V7GhYj0jhR0vT9aLMN9i6hhsvwNBQVAqK4JE4HK9vqk+XquoC9PbePhCFYVXf+YLf9TDpKOf0Q8F
CfhRR/VuJCXsXHYPE0JZrmzfIaMMNfWuAZSM70Xtst1HzQuUdCQbN1ZQBbfq8umt5oyBySCSVbXO
Mp7GfAx9yyaSo9sItrDpPM8hZarzoU7URY1+fj2BWnYJag9kwpUTB6VinWS51Aweh0EjeFd69g7E
Ujfo+B0rxLUDqPIKYg/7eKcfteeMd8CFou3t86nc5+cGqjH9OJbjGuQBqQcsfOFyqtx5HDDWTWqU
KbiTnOo2CJvuuE83YzCSnnFmQx+NA5lPg64+yTW06QJC+0Wf4SyuPy68kP7fIsYzoKGUG2M5D1+b
4PJ1G6PTrpaRAxGDLjvB5DDcPDWrXMnGbjSjNuikmbb/HPWucc22ZOCsabnsXQTlAVFHTceTqCC2
O5Fr9CZ6JZCYuiwiTWnQXUATZj1Lw14azl8UoPDrUwNXM6gSBsjWzVtbn7p4s0ADMRkat9zkzLjA
EcNvmUcjwnkP6DiXD3iBzdpbt+NoiZ2eUBLEiWpeVFmvROl9GBNitb3XY/cpqxqVPFnjp72cAWTT
kDDsXI4kAYA04ucAEG2rfyIzMew5/xU3/Av74uGeK/4L2e9QWCp7VJTSza2XXvdXbvjuaGA3rJVc
PPaAUgZ8Kb2OflYVqcuja1uMfUPffcqe5AvQd+w04OiLd42EnFFJk6CHlXOLwMZ51GKMVp7tMTkL
m8wTMJr32Il50Yipkwg/RlLyYe+C0CJGyBZiqK6/MkzMinj+3ph+Nh9Zd/szM0+EbyQRVgjePpng
sXKr9AM1RnTo3iEkLZQ2OsaGIPTDvulowkqkA9VwX9uOAz0B/tsCPICTT3PWashMP0x+CFCBpVHf
0EZy7RAbnNQW6WG5ZXAaUnx+dAlf9Y45kgcJJMP7YbiwwLev8pJid1PHI7qNFS8GJAvI3JLGvd5p
2S7GYT6m82pdKoOQhr8v0aR9vxYTVoAd0T3yp5e3mnVy7H1JVFsFgnvLLTgJFEf4f1Bu6Q/5I9ii
GZFssgxHt+JarhrmoK+NpwsTjcwsjUAre9oXhwOsy/6RX7jGGBeUNI3m+Ul5aYrA0Ju3uZV5mUeu
j32LYaO4TyjEp4eNCu8mrauasFvwNtDvsDH1xTcbi/Ch+uq7o7YPRQTxiUDpFRE5Nf75a/ZEHJDy
lTZ4mMuflyvxu8/xfd3OZpaJG2PB5hHRtyC9fK3CQ1NOHW8aYATbAtEX+dRjSbPHRP2SkZLCZosB
kRzOx++EcUTqvx4l/FLQj06hK6qJBOaqmknNEX22/Wslsi6fDKJCB8dKvNpQWEoSqz8DHjOJgTsV
4UQUveX4jF+d7gwwQXaHnNXV208POb5TdWVjgdABaKbLFPh1524GyT+EUrxg8HxdUN0kNctMCRz2
1niTwmHnXhlRXwMemEhYp0RjevZu/sirJj4AgVvYgC3IVuGJjH/ceHOWDAqtqFv6D6/txAhWokHV
uYlL8ANjW94GMpqTAY2Btqz6ar4ZrRsK5Xk7hvN7m7AvN2SXWFB1eUKTFCPnah9UWBZtnUNWsq8F
HvETCEGVu9twzPYg9LLase2ngHZ12apU3G4nENGl2VciD3DqY5mvfRL/kwy2zO13XwNOUgBhFVJY
bjiWQqz8XqQdCCOLzAmP7tw5octMdWinMQyX6BzVbmzWubMasrWGmrV2ziybI6YtEtnioQrIQcwZ
ZbNllXlg0Q7U3HDO+6rSAUGjNJLOduT6bVHKw9uhaq1mFbcjtyaWcrGccLrJopQaN2LqNFoGzELw
wxOlUCg9R3Qt8wPOUfkk/DWEOcd2JcfI5PkmdxCdP1l1gsxAlw4fg/iWM30iWf3YoaiGCB57yjIL
StB5of2Z3idM6CM2+mSA5z9Zrs7XW2WY3Y0hb+rtpV3c5fz6UpL/TEi9yXkr5pII14L7voBqCxuV
/EArsjmcxEtYqG5hSiQZ8+YOIoNmK011SqL3xu49xiGL7TrUqZQLM/Ax+I5kJJ89tnszQCHePg7b
1L58OiW+2enC0dAD9ECYX+BVvYBwx6ZMHj03FAdy9PRo7RDKd96j89oBCAIjVprymkdHRdgrfXfg
lcHRxlmGHCYrJPbB5gxVjxjYBSLTasmAj9VjtfHO5X1gzpWUGLkShcntl8aV41dM19HEgfqbo9p4
bmCyFXtLEfophLwzVzY6mkNZ0QNcaRLDE6QhSl2PLlsNDWUmANagl5UT6SsTOTL3f++CYvN00nB1
HDLm2ao+8zy9v9ibcS0bZJyxioqU5Ki5RcHm9LqAUs59KFDXCgXTGNxZFz5j6Ia/ZIRE99bFLZjF
AGwOS1xB10I4vbDW8Ina6SvR/1w0gIPF6g6v9TovsTMAszI9k91m7DUfdjgqlInVaSy7A+OGZI51
XcYN02d6N82cbnUeqQfPy9mCAL5KNm9jYCikNAkMZX+cxkaRp5CubaAZX5Hmy9s+9imOKU0HpvOY
MDxNxe+E8ZQXQDuCzc4j3WB8epbqPQtH05EorGdJPEcqXPcw/WGztqxJq/CUFuZU+3PoEOQPuqgh
x3lUfXf7Yf+ulfJFI/DNUWpT0EoCEfi4gS39q9C+DlXBdgYHauna6ugzi4FzQz9mNOZXB+ZSi1oY
q6C17ZKmo3HKe8nc1eKjq0QOl5xLUOkuQtvVXKwVZYhpWF/8QJm2KQFkLAoVCQXY35Bq+POVX60A
ZNF6HrZ5JYGAYQvxX4ed8Mge5GN/pYkjMAr6aeeFsZ/u1QZMBEzslvLEzaIRl3ftkneyoCx/41MA
fVCvVlRUUQxHByO8gTOIp7bdI+TK+Vz3zhvV9KM0mxxXgks9DVbIHjaiLNHnVKH43CdqbJ7m5KuC
gtCB5+lfpMfWoyl6nWk8VcAGJA9dHdH2JC29ZyywK8z7JMJl5ygI1aLmfi2Eomd25EMa2JszN59/
3ay45wNCjgKnnrnT3JYSy3rjZCCZqw1GWqD45Sqrva6/ovwQgj3oOTQDsGbAUHPKAz+3eAWd/x2B
Y15zlF1x2RUDtify2MMgUfsuj0DriCZ/j7ryqi8HW3iRBdq7slDjFzGbC5+4e7LqI92IAfN9iOYq
EeS278tngONW+9armzUI6vDKQz/i/uUqO4zn5u6kmIoXtYYSHK0dApZW6UF3gUDHm3KbmwOD1YLc
afg5pIOPiOf1Tdn+nt1CAL3sKu3J30GN+0xeCLD3FQs0tePiz8M2yRS7eqjKxXUG0DSz0+o+5kbq
whne4pTTH74yV0HNLzsj+KfJ3QnAp/zqKpfLpc1aozNKGIaKRxte3wdu3oB0z/vICemNjlAnG2/7
mkzKWZC9U39Mta672GJo029WX8sgTdAJohdzBl78a0UWbjHJ15YsRxkFKhVlYSUgPiCw7wVQGJSu
5svVO2s/twvlA/W9kF6WEHaJ+OgzRx87bXhwNdQFofjzq+Vtoh7Ey2L6YXZaeTRKGvp8jb+eSYo4
pjFJcrhIAPRM0zTbE7kndvnMwcxCzhr8AdyohpZ8wcwm+pPALQ9EDhbc2+nLJCyz1Q0Gb8eX/X2q
3wcfHJ3NHQ/PatrD96IqIxLFBzukejrhHX5HI2TZShvRbCPtDbPk57KqCOwWVl7JLDpypa7X+kwr
7raeN74pgJ1V84Io4yNEw2YUOOa4MO8AAVoymnnwdu5SCZGhSr08dWXUSqVOGvPxTRPulNStWRrM
XjL7BBSUgYo8w32mhEF/7cE+jgkuLnsXJoY9xXSEZh2/y8vsjzMJvbYilWBxplj9sGtKMB0AHF6D
tBib5Pup+pCYJ+24RE1SXytUyQFgnPfrn/3MhORbpnUL6Dv/gKvDSbSW3KXXb9Au7mBJ5O3HXJuX
azQ9/ghHV0rJyRtQE9Pd0RDwKHuqQzsTexMNOlQApampySc8Fa2FIeZgmSHzlmxKMRbZljwacYxE
x2gdW6yznSuuPAps7RdKxeMtZigDZRM0EPIY9RTM68GmqfVnx9fapWXQoRVucD0cRx1ku3Y6xU7Y
WqWOKcprzUFrajGdlQTZX4rbuh3lXEXbCAs3LdbeAGAsJBwr0ezTLs+BUKYRvF6u9dQ0vSiLoFrj
SK0br/TFnYBXcGCZbKgfpqtfgl+u6aV8VGzSpSCSEwafL7AAbyp4B/H5+Mhmna+hpzaBLZtIodc0
v3IU2Yz5tqiyOkRTh1pbdPTdc3yevrAlf58vjU9dvUWqNKkcDh3a5s+y1Wm/2UQQKQ6H3gRhm1Ku
LwAMR0OAchmS/uJO0BoQtFF8OA8J6DZI8Qur6PWArEP9eO1jGwMdadiXAmwooo83QWV3oiZKGGum
irOjA1MLnVF7i3WTiui5Kb/X5I4jOyVkIgiil1++MdvbXhed/KDfXR0sI1h2uUn1jeP5G6rt01lV
Snic+1z2zBHJHaBkt+oNom5aZU9P9WozkGV58cybPCOAjV1mbHhRzT9yUASLEsV60dbZlKKeT+hL
7/kAWy5r5I9K/OqSZf9y8FmZpciX3Toiz0x2J3Z5YyEC6vgEA3rMs3j4tmM2zUb07Kh41eV9yjRH
tmm6c85TRVAjcG3zG0RD3i+/NPvLmcI6ckSezlteeHXC/nfF3hIaWANpSWHw8AqQ2ZsxCDMxgOIN
Xrn0SCWTfKNRNwnP3E6rcqLIeZtz3ln9w1fBGL3pDqvoiv9+uIRTp1qJlBNYD4zWTxoUUNtO2Wtn
4k35Kx5a4ZEi33CD9SwLvj//s55zx1EUesKTDRR6wn6rY6xoKbmwX+N7t0WeKogsCMDael0hVSB5
iCO3fZ8xBBTDtWg87GdBHD1r6phk1HPEB9U1MwxjgU/656I25zYeALVReM8alUbeGEZPow5DBkyr
Rs88iiXx3ra9D1wDkqBm2eOcOp16YUwwbXBbJgjDyxwBwxMV/B2QW1IbAaWWkpKFrDuA9Nof43B8
dPnczHymscny7JHQz2YKWGYnHNjb22t9zvsBcizNlOazulgiN1BC4rHSPSbjU49Ec2e2HzGuAuyU
0oc19K0a/nw900qxnpeNinPazxUz+lXde6lGiaaRiWgM0xrPL7+mdhb9F/jx8wv0pGSrndRblttp
TVNVlQGTXwi7JMLaCmZBIeIEEbrIJgmRzs7uh0HmMrgTBKu6Qsiqvp/12Vl6RETh1w2iTFTwt4nT
5h5n520h3jm6meFOw2tp0n3sM9QdzJ7mv7b2CgZiG8r0WkCBfCyXBpQu9igybnFrO+QJcREAOY/h
cN3mz2y6xbwq2+9TScwe9nPTec+bQCezmGFfOnQtK55gnhNLof9y9K8cK5NM1Ttsq2QL3xbsQg4p
tGipN75CIVQ1taU1kmOnmIWjraODL0F8tmbOX9GotnNf0GcGA65dM+lYu3TVM52wVcujmZeKqAgS
4FEShW4TUS6Qe3kYq7khwKv+3sIPof5rp2VJnVSqGI6bbLPHPugmTLertvmbl4pSDqCcj4OfX6EY
FlkaXtBQUFRGgJnLpLqVG6c7LW/di4PA/M4StkJIij/j2huVwXNQ86zqnV4VflZUQCIyFGcGY3B7
LOI3EBcVhOTYmRY8Y/SAdQN9fkbQJkIViwxfDAM0iSNTz48PJDTO8kqOGAP9R2V6mtP6sqJWtLz4
BKwlA4SYF1/dfOAWw7Zt+i0lqOJjRiEEGH4iYmR4QYEVhMdOvgUbqRYB4S73xdRIUQZlXAxK/eIR
R1HgtqNY733yCkjDkaZsHSDIimecny83UvLfAavuamXjsdSPOiLXdCoRp7I1wbeA/yIYjZFATsE5
A5oJ2NZJSIhUzBLtbYwmzfk0hW6uY0/1jfOPpN1YI/wKAPSmaHtUFTqcTGQ905ih/zQmBaRF/pyT
AFV6s6PecrHg0T9M602Dd9Ts8Oszvtaa73pw84dC/OA6RaPXj7GTpUaXT28GY7fFwOS5oFo/aP78
+mVhhE6Uza7BNUcRPFms1RtBm/Y7lC8aGnMu5cA5qWcM/nrE3j0jonXFiZ78U4MyhtFCGk60mnpx
AF7jD6anM5r3CZrWSYs4bMfQA3FO34kau70EZJEkMSbwEGLgnRDKc7jN/gTUMJ/NCOMTivTw671N
GPuOmnzxQvFrmtFIfKWEz1XMfGKYoqj9E1KVAoMJCDOVw3lzjbsXq8EHlOUYhSo9pDQwCJsGDyy8
j1CVVz8a1Cn3F6LvOsBpbopLa3Qfx2T1M4NPd/CJRXUrFTenfr2dL5C8eImA/czrO2p0Gupbjdyw
ra5K/BjCAqHjamOTteNEqfwNg/GY1D6bnWUW6er+9kBPJsOBffbz3mmbpWQ+7AslvmpTVDa4XA6x
+lMpXUu1OPEwmC1/HjXWycgT6RheZi2Xva/i/xbQSffnzX6iqWexI72oj9FEFfzrjpKeElefdLw7
yPIsO2AW4Tx4Org0QwA4uqy92VCq/9T2em1Gjw1RSPYy7DpfyB/hgcBW8ga/8pXIZwSKgcyTlFKT
na/ofVjs7hmDlBDkizHely6kYF+Xp0L0fZFohwjGPrIGfuD/FX1aYI+Gg8rgBv+FL4JXPnveTyfw
2slPag9Ke8Htdfh33FaAhhcAmIkNri+v5kvEoKncf98Tcdf7Gmn1IGjPAd2Y5U8Exmen9ylYtqvy
7mmK2K+Xdm+IzZCjEp7sMUPr1Ts5K+zjcymF3tfKj/DNDx7ol0tFIZ8oVGTvoIlXa44ntzYCstZ1
uzXLgKU7uztio07QPX6EOAMLzILIG6pQy3ISEE9Wonf89iW6Arg5K9HfnsHIIFKSuqCGxidX/Ef0
ywFocbUyWl2T9e5VIxakyjbYS1R26mAZO2OpITr9BuG3QXDCD9n4Fi2pTPg3GPMEjvKz82jC3+4W
StiLs7M1A5AsFhcxOC3q4wQ0AFScmRKOpCorTI8aa8xm3xTjF+e6kmux14X79FK/0tV1Tb4yirwq
j0CpKLHIp/ADoNlF5gqpp4wIhGTikcjHxhfBlAuSUnw1opSM2h5y1eU7wmvOFhzvQRSraY79Y9vQ
s7HJCjgMPZKZUSNb5UfBufgUcOukBjI9OxOU3oc5cMNXrSApVH/rDSKYg7ZZDu3+brQJT2hTeEcL
meyU9aNHlaedP8OtDqQXaAIN7DtD+SNHMk3AlJTMNt3ywzx8WTuKm18ftqRp9j6Ox6Lwr3XaRPXh
gnjZdHaSbrt+Mn/W6lHCAyEBKFDPQWOfQlvojIjk50L60HpMmbPS4iQhBeuxJK3+YDisOUtshhGZ
C4iuugNosJDogL7/D5YTSbmYYqOWOLddWuDTReWCweuWphj9n83Fih7wLh5lvOim7rJplLEHrcvq
0PjHwRjF5Fev5OynNW+7N51DIRwVNDjyRMGzXAutHxl3cCeB5ccTIGxKCnlG2vuPt4RCes4La5+V
IsHpPPLxrYSPjUmLJh+qBZKiqiI+sM83WcASdRbBw8HURXGaPQf/zjJz3SVQxmTFqweCGA3bw12M
Ux2ojHAljlN3awDP+oLRugvnUdg7vUsZ2aBDECJag358bzR1vwlrDccE+7KMno+ZJ4A3ED2Vqs3K
Lv/84lK5v6mcJHGbzGpKhNo3zHh8IyluAhfn1ZhTgvNdBL+SzmOyNQoK8/5QaaYwvi8Kg/Q+pC+j
Z+qjos9wMLVwnUpDlblAVO0xRzWkdMaCcEvJhBPZkFZ1zoLEQF43u4vHelODCIO53x+aNo1yV4Eh
p4dKi/Zj4vQ7RdiC7Qbb3Lnf+6cZznOYeKFsy+kQF1MbP6sqvOqgB3mv3exp078MX7W9SrJLYjjw
baudlfj+kKBYj5OPazOpTHBwVL8Sc+D9OIj4Wko9QDBiKmaZNLJNmUMNBHScqCQF6mepZX1IzsUr
rFZ+faXusIZflxaqvo6XsLx65b67NPxT4RJXO/nsfsJSuDeQjhSg+PNX0mRXiX47QYQvR6xLH3i3
NPoqDR3EFGVNKgfcXrMvgjSfPMdn3CZJF8Z3IIB6ZNiWjudNbN5VQZ5kxJGGFQk1qeVuKU0EojhI
CRqExBC+y0So1ZFolTRiFz9uu1q3Kr1Hu3xMkW+PcBTV+4ZeeMARwcKRqcQj1gnfQZzQBnYsWcRN
DjKU/jpfwVOiTBb7sfDlL3XVSCqED9hkSgVa7sZxR+Eyel9wWh7SmKroqiTEJaX/th8qDSUzeBcO
W3ywg/OlB4+WPs8kx44xsZQtRtXfGQUUt5pDnZFHawdu1ULzSvK4lkRjlGEyXO+B06D44KMcd2J7
Vmi6R5lhkdg3/7FpjEZhOYqKregA113SY7WkmSGi9AJ5kXZepeONPuv7CZontCySr1szzEeNS7yG
WBhr29Wpl00HnfGyWK2FAxld6Q7i8fk6gSNHCGdwGq8pOBE/+XO0UyBf3DruN9gCQAyqNxn3un0w
4+uCCDsqO09pyFdNJbZ5uwK4flTDQ42JpllZQXxPJtxR0H65fWsBdu8tgRqO8a0Amx+GUxf0dIew
pwO/s2cRlpQclaNOjjGZ1YQEshx/Jt9tPFUVkDQc1kit9Y9MdZmhSJ8HROVRwbW8zC+XrOhrNrwc
rMz25wG50tG2c9Wu4wJBFKJWHwalUpsMZatbOaFrp7p8s4jlgAvi0YBEyVG8H458OH1Sw5gR/zax
5bfJTrzJUNpyzm5nL5JFR29I5HktFUpekmsEP4z6qL3U+BCJQbhs74ozL1bfwOmR++FWvhHW+bys
AT+p5CUWzkyzPoxADPzgtlyH9RAuI8SaRCQYCXaMgofvCSSXqTMJKxXP6r9sdbC9Yp9Jif/N1KPX
nSBycHrqnPAh8I7nW03qWbt83QMXV6hprEtP2ZhSnA9zpvq3PzETo/jVakZDzSf2SPYlish2qzJI
35vq6SixVTWj/MgLz1qSkkoAeb2zmjeqHc0Y25QSHbfqz0APa7eDVdT/G/j2X7799NT17w8Vc0Kl
PpIi4OpIzwTzf46hsRRvib2FRy8d/QAXI3L04/25VxDRTsS92vI8bK9bz/CjCa/5QkSceJLYUwu9
FdFUzUmiDJZRRBJoinpYwkLXCo7tm2PXbm9g7QfsN/zqsHkUCtikV89ueyAsCKCGeMAkE6Xz3BGY
4sU1MJAVPwmKv/U9gEJD9ji04Zd5gHQq/Mn6corm1MbO9M9qVFfuenWMqeogJUvhGH3t1h2FcfWe
gfrDARblfbOyBoYW1QLT8ybHQQp1MWfBVbSt+vMuyCzd6DwkFBObyToj4KhuNmTF1JlQh/0/QsJh
0JPLMkw3tKUNROhudby6vALHpzd5r8yRnlFTDG4SH8kXFoDM+VQTFGMRxu4Nsiov8bRC9S9wi/ZG
Wm5ODAKuCSQ4JTjdyDQYFS0gP4SswSxlxqYnr4SaHCpRq/v4MAY80GQsGxLtwggqSohwhq8n02oo
Y4gsH+HypWkiC0g7Pgfcq3xYzR9WcUTzZu8QH42kSSBcLTRLiCD19uH9wfxNNsW0Q9rs+UodGTqM
iyZzaPA9g/jIdAhBkJ5CzUyOVlHcQ+SgGR7aA7q7/lBNhvYvSH4AY1blY2v3qXH0zH1V6cnKJddh
QYjZlZtxvVF30EityNNNcwRyaYuwNKcJs4CzHwOmlwv98Q8E+FekW/Up7T7Zlgdwtq32OxmDPkr9
NXC81vbf+kUsujW0lYaKhK1fHc1LDFwlKcoauLaKMwVfGsEJ8KL6v9Toixpc1tIz9LgVLPERVwSs
qIzNq4BWe4pvykFhPXS67ul9D9+HgebWtnnKCuMoTszsG0aNHcgqTrvm6tnqTVV63CqZZr1iug/H
+CIcNEZpmqC3XSaGSemchwzNCBCPLJpsPLI8s7KulHzfpGDAjiRSn2GuPlhxjT8CTcjUD30683i+
fca14Jed+SfeL4QnFlDYtBAIcS7Cwd/cPzIgsU7GTGM8WVgsDaUpfXWhTzBtEhOMhFZ2UHa++X08
ooMFbLPyq6t2nhSE/eJZg4cGWcyzwp/ScNRf1Yi2QBwIUO8Bfe44/NKjoklyj3Mk3ePwe0Iv8qVC
4WcY00HZMqts8T5khk2yzCAlkItOr03Afxp7e3wIH8sAwlmrKbnED5+3ANkbLAe021f4+pPLlnHn
lPSwuWKUqJOZbxM5g4GXDJCQ6kobqPSRj2UUwDnLkbf44sVocPLebURulC6Nf1NNY3sG14XSxbP2
j2QF5XsHV4dWHFJ77rqERc6LJa7Mq2UHTFmI2Lev6/DvVsjyytDktJU2XmA3O+U3t83TzTFBsnhI
aGZIMT5eeaINas4xYW2kPQCdxPm5fbW2bZocjr2M3QPuCZADZJuP4m0dKbK9gIW57ACFzZ4U6XIA
Vf7fFMl2ic4cazx4uA28RVevEVI3Nq8+aZHIxe/1jImhj+I2UWXzPgKwh63zAPJFIP/1ACHQaNBh
8/EOhrmx7ca3hdNI2VbLpm4taCJ2KMhnTNAL7bvl+ckXcf9+nKiqbSglTPVLPNIAGBXiV4VUnovu
IALj0f/cXCb7xJqDdRTLV4FAbZ+ldO4m3riv3C1SbGQTu41PCk2m6o1OEoJvqRbCWo9T4NGQrgzO
wqekZjXCq4w45DQIZZPGGwtgcqvEzy0P/hXmnzZw4tsabsmIKaiT64ip8T6kjqWpadgyNMnxY4vJ
W5KOYv74i9+eKI6PQKvkSTWgECxnnTHqMmY4JjGpMAQ7MHdWFf3b0Hunq+SmBTJFQsS2EzzUAZaL
bx23F1e6hIK6Gcbx/6itGfZEamphcXBYgM7zpFDe4kdci3PghD+WyMa7c3i5+x+f0MW8eQhBXqKq
dZgKYo7EP3D/46OX4goHi6xZD1/LACL7CI8UuOilb3296S4rHwuw/PHgBLm0GmVfLOQ0s2mADqEM
WSY+hYQGwtHsyHaLfGbcYqf2BPpcXNtpdRXAE/LxDpJzn5hbLquwVuokLFZJjQDVT8Pce8HRP0Y6
gl/K8ud08Pw9a/5u+sIjzTirMGRypD1Gtgij/lTWpqok8HPVOgNwEB5TvBEzvDGWMj+ZcA4EXo+Q
iE7Rqt5CLtfD9Z7gOcGlZW1s4hFkPaEZ79xxTuaDWaxHCxpBaDJiCnWAnFDf1j0DR267mAP/tbK2
JCfTE54bo7moS+cVpYJS0FuwBEDqs/SZpbkGa2oRGk8btfsgVNlgYvalWXujnK0f0kEauymaPFWz
4jnGGZQbwEbFLZ+LDoNPcwv4DdvjjAyFNnmvAvbwQ+P2MV5TfgYTsbpdPqMyhg==
`protect end_protected
